
* Circuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 ;CMOSNuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 
* TDB File:  C:\Documents and Settings\Owner\Desktop\Project\Multiplier.tdb
* Cell:  Cell0	Version 1.10
* Extract Definition File:  ..\extract\mhp_n05.ext
* Extract Date and Time:  01/30/2023 - 20:29

* Tech: AMI_C5N
* LOT: T22Y_TT (typical)                  WAF: 3104
* Temperature_parameters=Optimized 
.MODEL CMOSN NMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6696061
+K1      = 0.8351612      K2      = -0.0839158     K3      = 23.1023856
+K3B     = -7.6841108     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.9047241      DVT1    = 0.4302695      DVT2    = -0.134857
+U0      = 458.439679     UA      = 1E-13          UB      = 1.485499E-18
+UC      = 1.629939E-11   VSAT    = 1.643993E5     A0      = 0.6103537
+AGS     = 0.1194608      B0      = 2.674756E-6    B1      = 5E-6
+KETA    = -2.640681E-3   A1      = 8.219585E-5    A2      = 0.3564792
+RDSW    = 1.387108E3     PRWG    = 0.0299916      PRWB    = 0.0363981
+WR      = 1              WINT    = 2.472348E-7    LINT    = 3.597605E-8
+XL      = 0              XW      = 0              DWG     = -1.287163E-8
+DWB     = 5.306586E-8    VOFF    = 0              NFACTOR = 0.8365585
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.0246738      ETAB    = -1.406123E-3
+DSUB    = 0.2543458      PCLM    = 2.5945188      PDIBLC1 = -0.4282336
+PDIBLC2 = 2.311743E-3    PDIBLCB = -0.0272914     DROUT   = 0.7283566
+PSCBE1  = 5.598623E8     PSCBE2  = 5.461645E-5    PVAG    = 0
+DELTA   = 0.01           RSH     = 81.8           MOBMOD  = 1
+PRT     = 8.621          UTE     = -1             KT1     = -0.2501
+KT1L    = -2.58E-9       KT2     = 0              UA1     = 5.4E-10
+UB1     = -4.8E-19       UC1     = -7.5E-11       AT      = 1E5
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2E-10          CGSO    = 2E-10          CGBO    = 1E-9
+CJ      = 4.197772E-4    PB      = 0.99           MJ      = 0.4515044
+CJSW    = 3.242724E-10   PBSW    = 0.1            MJSW    = 0.1153991
+CJSWG   = 1.64E-10       PBSWG   = 0.1            MJSWG   = 0.1153991
+CF      = 0              PVTH0   = 0.0585501      PRDSW   = 133.285505
+PK2     = -0.0299638     WKETA   = -0.0248758     LKETA   = 1.173187E-3
+AF      = 1              KF      = 0)
*
.MODEL CMOSP PMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9214347
+K1      = 0.5553722      K2      = 8.763328E-3    K3      = 6.3063558
+K3B     = -0.6487362     W0      = 1.280703E-8    NLX     = 2.593997E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.5131165      DVT1    = 0.5480536      DVT2    = -0.1186489
+U0      = 212.0166131    UA      = 2.807115E-9    UB      = 1E-21
+UC      = -5.82128E-11   VSAT    = 1.713601E5     A0      = 0.8430019
+AGS     = 0.1328608      B0      = 7.117912E-7    B1      = 5E-6
+KETA    = -3.674859E-3   A1      = 4.77502E-5     A2      = 0.3
+RDSW    = 2.837206E3     PRWG    = -0.0363908     PRWB    = -1.016722E-5
+WR      = 1              WINT    = 2.838038E-7    LINT    = 5.528807E-8
+XL      = 0              XW      = 0              DWG     = -1.606385E-8
+DWB     = 2.266386E-8    VOFF    = -0.0558512     NFACTOR = 0.9342488
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.3251882      ETAB    = -0.0580325
+DSUB    = 1              PCLM    = 2.2409567      PDIBLC1 = 0.0411445
+PDIBLC2 = 3.355575E-3    PDIBLCB = -0.0551797     DROUT   = 0.2036901
+PSCBE1  = 6.44809E9      PSCBE2  = 6.300848E-10   PVAG    = 0
+DELTA   = 0.01           RSH     = 101.6          MOBMOD  = 1
+PRT     = 59.494         UTE     = -1             KT1     = -0.2942
+KT1L    = 1.68E-9        KT2     = 0              UA1     = 4.5E-9
+UB1     = -6.3E-18       UC1     = -1E-10         AT      = 1E3
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.9E-10        CGSO    = 2.9E-10        CGBO    = 1E-9
+CJ      = 7.235528E-4    PB      = 0.9527355      MJ      = 0.4955293
+CJSW    = 2.692786E-10   PBSW    = 0.99           MJSW    = 0.2958392
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.2958392
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 5.292165E-3    LKETA   = -4.205905E-3 
+AF      = 1              KF      = 0)
*

* Warning:  Layers with Unassigned FRINGE Capacitance.
*   <Pad Comment>

* NODE NAME ALIASES
*       1 = U291/U240/VDD (706.5 , 307.5)
*       1 = U291/U239/VDD (681.5 , 306.5)
*       3 = U290/U240/VDD (422 , 307.5)
*       3 = U290/U239/VDD (397 , 306.5)
*       4 = U290/U240/vout (429 , 287)
*       4 = U285/U238/A (872.5 , 224.5)
*       4 = U285/AA (872.5 , 228.5)
*       7 = U289/U239/VDD (113 , 306.5)
*       7 = U289/U240/VDD (138 , 307.5)
*       9 = U298/U234/INPUTA (-1067 , 275)
*       9 = U298/X (-1072 , 289)
*       9 = X0 (-1072.5 , 287)
*       9 = U287/U239/A (-758.5 , 284)
*       9 = U287/X (-764.5 , 289)
*       9 = U293/U234/INPUTA (-505.5 , 276)
*       9 = U293/X (-510.5 , 289.5)
*       9 = U288/U239/A (-177 , 285)
*       9 = U288/X (-183 , 290)
*       9 = U289/U239/A (107.5 , 285)
*       9 = U289/X (101.5 , 290)
*       9 = U290/U239/A (391.5 , 285)
*       9 = U290/X (385.5 , 290)
*       9 = U291/U239/A (676 , 285)
*       9 = U291/X (670 , 290)
*       10 = U288/U240/VDD (-146.5 , 307.5)
*       10 = U288/U239/VDD (-171.5 , 306.5)
*       14 = U293/U238/B (-371 , 300.5)
*       14 = U293/U237/vout (-385.5 , 284)
*       16 = U293/U237/Vdd (-404.5 , 307.5)
*       16 = U293/U234/VDD (-431.5 , 306.5)
*       16 = U293/U238/VDD (-309.5 , 304)
*       16 = U293/U238/A (-277.5 , 302.5)
*       16 = U293/AA (-277.5 , 306.5)
*       17 = U293/U237/vin (-414 , 285)
*       17 = U293/U234/OUTPUT (-425 , 293.5)
*       22 = U298/U234/VDD (-993 , 305.5)
*       22 = U298/U232/VDD (-906.9 , 303.1)
*       22 = U298/U232/A (-874.9 , 301.6)
*       22 = U298/AA (-875 , 306.5)
*       22 = U287/U240/VDD (-728 , 306.5)
*       22 = U287/U239/VDD (-753 , 305.5)
*       28 = U285/U237/vout (764.5 , 206)
*       28 = U285/U238/B (779 , 222.5)
*       29 = U285/U238/S (771 , 223)
*       29 = U285/Sum (771 , 192)
*       29 = P1 (915.5 , 185)
*       31 = U291/U240/GND (720.5 , 272.5)
*       31 = U291/U239/GND (711 , 272.5)
*       31 = U290/U240/GND (436 , 272.5)
*       31 = U290/U239/GND (426.5 , 272.5)
*       31 = U289/U240/GND (152 , 272.5)
*       31 = U289/U239/GND (142.5 , 272.5)
*       31 = U288/U240/GND (-132.5 , 272.5)
*       31 = U288/U239/GND (-142 , 272.5)
*       31 = U287/U240/GND (-714 , 271.5)
*       31 = U287/U239/GND (-723.5 , 271.5)
*       31 = U283/U234/GND (100.5 , 194)
*       31 = U282/U234/GND (-184 , 194)
*       31 = U293/U234/GND (-481 , 272)
*       31 = U251/U215/GND (894.5 , 73.5)
*       31 = U251/U211/GND (792.5 , 74.5)
*       31 = U249/U211/GND (508 , 74.5)
*       31 = U249/U229/GND (421 , 124.5)
*       31 = U247/U211/GND (224 , 74.5)
*       31 = U245/U211/GND (-60.5 , 74.5)
*       31 = U279/U211/GND (-345 , 170.5)
*       31 = U243/U211/GND (-345 , 74.5)
*       31 = U279/U228/GND (-481 , 169)
*       31 = U241/U211/GND (-629.5 , 74.5)
*       31 = U252/U211/GND (792.5 , -21.5)
*       31 = U249/U215/GND (610 , 73.5)
*       31 = U250/U211/GND (508 , -21.5)
*       31 = U250/U229/GND (421 , 28.5)
*       31 = U247/U215/GND (326 , 73.5)
*       31 = U248/U215/GND (326 , -22.5)
*       31 = U248/U211/GND (224 , -21.5)
*       31 = U247/U228/GND (88 , 73)
*       31 = U245/U215/GND (41.5 , 73.5)
*       31 = U245/U228/GND (-196.5 , 73)
*       31 = U243/U215/GND (-243 , 73.5)
*       31 = U244/U211/GND (-345 , -21.5)
*       31 = U243/U228/GND (-481 , 73)
*       31 = U241/U215/GND (-527.5 , 73.5)
*       31 = U242/U211/GND (-629.5 , -21.5)
*       31 = U294/U211/GND (783 , -117.5)
*       31 = U295/U211/GND (498.5 , -117.5)
*       31 = U297/U215/GND (316.5 , -118.5)
*       31 = U297/U211/GND (214.5 , -117.5)
*       31 = U310/U211/GND (-639 , -117.5)
*       31 = U302/U238/GND (-880 , -91.5)
*       31 = U302/U237/GND (-967.5 , -92)
*       31 = U269/GND (783 , -168.5)
*       31 = U296/U211/GND (498.5 , -219.5)
*       31 = U296/U210/GND (498.5 , -168.5)
*       31 = U307/U215/GND (316.5 , -220.5)
*       31 = U307/U211/GND (214.5 , -219.5)
*       31 = U307/U210/GND (214.5 , -168.5)
*       31 = U304/U211/GND (-639 , -219.5)
*       31 = U304/U210/GND (-639 , -168.5)
*       31 = U303/U211/GND (-936.5 , -219.5)
*       31 = U303/U210/GND (-936.5 , -168.5)
*       31 = U303/U213/GND (-817.5 , -169)
*       31 = U303/U215/GND (-834.5 , -220.5)
*       31 = U304/U213/GND (-520 , -169)
*       31 = U304/U215/GND (-537 , -220.5)
*       31 = U305/U210/GND (-354.5 , -168.5)
*       31 = U305/U211/GND (-354.5 , -219.5)
*       31 = U305/U213/GND (-235.5 , -169)
*       31 = U305/U215/GND (-252.5 , -220.5)
*       31 = U306/U210/GND (-70 , -168.5)
*       31 = U306/U211/GND (-70 , -219.5)
*       31 = U306/U215/GND (32 , -220.5)
*       31 = U306/U213/GND (49 , -169)
*       31 = U307/U213/GND (333.5 , -169)
*       31 = U296/U213/GND (617.5 , -169)
*       31 = U296/U215/GND (600.5 , -220.5)
*       31 = U302/U234/GND (-1042.5 , -93)
*       31 = U310/U228/GND (-765.5 , -68)
*       31 = U310/U210/GND (-639 , -66.5)
*       31 = U310/U213/GND (-520 , -67)
*       31 = U309/U228/GND (-481 , -68)
*       31 = U310/U215/GND (-537 , -118.5)
*       31 = U309/U210/GND (-354.5 , -66.5)
*       31 = U309/U211/GND (-354.5 , -117.5)
*       31 = U309/U213/GND (-235.5 , -67)
*       31 = U308/U228/GND (-196.5 , -68)
*       31 = U309/U215/GND (-252.5 , -118.5)
*       31 = U308/U210/GND (-70 , -66.5)
*       31 = U308/U211/GND (-70 , -117.5)
*       31 = U308/U215/GND (32 , -118.5)
*       31 = U308/U213/GND (49 , -67)
*       31 = U297/U228/GND (88 , -68)
*       31 = U297/U210/GND (214.5 , -66.5)
*       31 = U297/U213/GND (333.5 , -67)
*       31 = U295/U228/GND (372 , -68)
*       31 = U295/U210/GND (498.5 , -66.5)
*       31 = U295/U213/GND (617.5 , -67)
*       31 = U295/U215/GND (600.5 , -118.5)
*       31 = U294/U228/GND (656.5 , -68)
*       31 = U294/U210/GND (783 , -66.5)
*       31 = U294/U213/GND (902 , -67)
*       31 = U294/U215/GND (885 , -118.5)
*       31 = U301/U234/GND (-1042.5 , 2)
*       31 = U301/U232/GND (-915.9 , 3.6)
*       31 = U241/U228/GND (-765.5 , 73)
*       31 = U242/U228/GND (-765.5 , -23)
*       31 = U242/U229/GND (-716.5 , 28.5)
*       31 = U242/U210/GND (-629.5 , 29.5)
*       31 = U242/U213/GND (-510.5 , 29)
*       31 = U244/U228/GND (-481 , -23)
*       31 = U242/U215/GND (-527.5 , -22.5)
*       31 = U244/U229/GND (-432 , 28.5)
*       31 = U244/U210/GND (-345 , 29.5)
*       31 = U244/U213/GND (-226 , 29)
*       31 = U246/U228/GND (-196.5 , -23)
*       31 = U244/U215/GND (-243 , -22.5)
*       31 = U246/U229/GND (-147.5 , 28.5)
*       31 = U246/U210/GND (-60.5 , 29.5)
*       31 = U246/U211/GND (-60.5 , -21.5)
*       31 = U246/U213/GND (58.5 , 29)
*       31 = U248/U228/GND (88 , -23)
*       31 = U246/U215/GND (41.5 , -22.5)
*       31 = U248/U229/GND (137 , 28.5)
*       31 = U248/U210/GND (224 , 29.5)
*       31 = U250/U228/GND (372 , -23)
*       31 = U249/U228/GND (372 , 73)
*       31 = U248/U213/GND (343 , 29)
*       31 = U250/U210/GND (508 , 29.5)
*       31 = U250/U215/GND (610 , -22.5)
*       31 = U251/U228/GND (656.5 , 73)
*       31 = U252/U228/GND (656.5 , -23)
*       31 = U252/U229/GND (705.5 , 28.5)
*       31 = U250/U213/GND (627 , 29)
*       31 = U252/U210/GND (792.5 , 29.5)
*       31 = U252/U213/GND (911.5 , 29)
*       31 = U252/U215/GND (894.5 , -22.5)
*       31 = U300/U234/GND (-1042.5 , 98)
*       31 = U300/U232/GND (-915.9 , 99.6)
*       31 = U241/U229/GND (-716.5 , 124.5)
*       31 = U241/U210/GND (-629.5 , 125.5)
*       31 = U241/U213/GND (-510.5 , 125)
*       31 = U243/U229/GND (-432 , 124.5)
*       31 = U243/U210/GND (-345 , 125.5)
*       31 = U243/U213/GND (-226 , 125)
*       31 = U279/U215/GND (-243 , 169.5)
*       31 = U245/U229/GND (-147.5 , 124.5)
*       31 = U245/U210/GND (-60.5 , 125.5)
*       31 = U245/U213/GND (58.5 , 125)
*       31 = U247/U229/GND (137 , 124.5)
*       31 = U247/U210/GND (224 , 125.5)
*       31 = U247/U213/GND (343 , 125)
*       31 = U249/U210/GND (508 , 125.5)
*       31 = U251/U229/GND (705.5 , 124.5)
*       31 = U249/U213/GND (627 , 125)
*       31 = U251/U210/GND (792.5 , 125.5)
*       31 = U251/U213/GND (911.5 , 125)
*       31 = U298/U234/GND (-1042.5 , 271)
*       31 = U299/U234/GND (-1042.5 , 193)
*       31 = U299/U232/GND (-915.9 , 194.6)
*       31 = U298/U232/GND (-915.9 , 272.6)
*       31 = U281/U237/GND (-690.5 , 194)
*       31 = U281/U234/GND (-765.5 , 193)
*       31 = U281/U238/GND (-603 , 194.5)
*       31 = U279/U229/GND (-432 , 220.5)
*       31 = U293/U237/GND (-406 , 273)
*       31 = U293/U238/GND (-318.5 , 273.5)
*       31 = U279/U210/GND (-345 , 221.5)
*       31 = U279/U213/GND (-226 , 221)
*       31 = U282/U237/GND (-109 , 195)
*       31 = U282/U238/GND (-21.5 , 195.5)
*       31 = U283/U237/GND (175.5 , 195)
*       31 = U283/U238/GND (263 , 195.5)
*       31 = U284/U234/GND (384.5 , 194)
*       31 = U284/U237/GND (459.5 , 195)
*       31 = U284/U238/GND (547 , 195.5)
*       31 = U285/U234/GND (669 , 194)
*       31 = U285/U237/GND (744 , 195)
*       31 = U285/U238/GND (831.5 , 195.5)
*       32 = U285/U234/VDD (718.5 , 228.5)
*       32 = U285/U237/Vdd (745.5 , 229.5)
*       32 = U285/U238/VDD (840.5 , 226)
*       33 = U291/U239/B (702.5 , 285)
*       33 = U291/Y (702 , 309)
*       33 = Y0 (702 , 309)
*       33 = U294/U228/INPUTB (687.5 , -62)
*       33 = U252/U228/INPUTB (687.5 , -17)
*       33 = U252/Y (689 , 63.5)
*       33 = U251/U228/INPUTB (687.5 , 79)
*       33 = U251/Y (689 , 159.5)
*       33 = U285/U234/INPUTB (700 , 200)
*       33 = U285/Y (702 , 229)
*       34 = U291/U239/OUT (689.5 , 273.5)
*       34 = U291/U240/vin (728 , 285.5)
*       35 = U285/U234/OUTPUT (725 , 215.5)
*       35 = U285/U237/vin (736 , 207)
*       36 = P0 (915.5 , 244)
*       36 = U291/U240/vout (713.5 , 287)
*       43 = U284/U237/vout (480 , 206)
*       43 = U284/U238/B (494.5 , 222.5)
*       44 = U284/U238/S (486.5 , 223)
*       44 = U284/Sum (486.5 , 192)
*       44 = U251/CC (759 , 161)
*       44 = U251/U211/A (833.5 , 103.5)
*       45 = U284/U237/Vdd (461 , 229.5)
*       45 = U284/U234/VDD (434 , 228.5)
*       45 = U284/U238/VDD (556 , 226)
*       46 = U290/U239/B (418 , 285)
*       46 = U290/Y (417.5 , 309)
*       46 = Y1 (417.5 , 309)
*       46 = U295/U228/INPUTB (403 , -62)
*       46 = U250/U228/INPUTB (403 , -17)
*       46 = U250/Y (404.5 , 63.5)
*       46 = U249/U228/INPUTB (403 , 79)
*       46 = U249/Y (404.5 , 159.5)
*       46 = U284/U234/INPUTB (415.5 , 200)
*       46 = U284/Y (417.5 , 229)
*       47 = U290/U239/OUT (405 , 273.5)
*       47 = U290/U240/vin (443.5 , 285.5)
*       48 = U284/U237/vin (451.5 , 207)
*       48 = U284/U234/OUTPUT (440.5 , 215.5)
*       55 = U283/U237/vout (196 , 206)
*       55 = U283/U238/B (210.5 , 222.5)
*       56 = U284/U238/A (588 , 224.5)
*       56 = U284/AA (588 , 228.5)
*       56 = U289/U240/vout (145 , 287)
*       57 = U283/U238/S (202.5 , 223)
*       57 = U283/Sum (202.5 , 192)
*       57 = U249/CC (474.5 , 161)
*       57 = U249/U211/A (549 , 103.5)
*       59 = U283/U237/Vdd (177 , 229.5)
*       59 = U283/U234/VDD (150 , 228.5)
*       59 = U283/U238/VDD (272 , 226)
*       60 = U297/U228/INPUTB (119 , -62)
*       60 = U248/U228/INPUTB (119 , -17)
*       60 = U248/Y (120.5 , 63.5)
*       60 = U247/U228/INPUTB (119 , 79)
*       60 = U247/Y (120.5 , 159.5)
*       60 = U283/U234/INPUTB (131.5 , 200)
*       60 = U283/Y (133.5 , 229)
*       60 = U289/U239/B (134 , 285)
*       60 = U289/Y (133.5 , 309)
*       60 = Y2 (133.5 , 309)
*       61 = U289/U239/OUT (121 , 273.5)
*       61 = U289/U240/vin (159.5 , 285.5)
*       62 = U283/U237/vin (167.5 , 207)
*       62 = U283/U234/OUTPUT (156.5 , 215.5)
*       68 = U288/U240/vin (-125 , 285.5)
*       68 = U288/U239/OUT (-163.5 , 273.5)
*       69 = U288/U239/B (-150.5 , 285)
*       69 = U288/Y (-151 , 309)
*       69 = Y3 (-151 , 309)
*       69 = U308/U228/INPUTB (-165.5 , -62)
*       69 = U246/U228/INPUTB (-165.5 , -17)
*       69 = U246/Y (-164 , 63.5)
*       69 = U245/U228/INPUTB (-165.5 , 79)
*       69 = U245/Y (-164 , 159.5)
*       69 = U282/U234/INPUTB (-153 , 200)
*       69 = U282/Y (-151 , 229)
*       70 = U282/U237/vout (-88.5 , 206)
*       70 = U282/U238/B (-74 , 222.5)
*       71 = U283/U238/A (304 , 224.5)
*       71 = U283/AA (304 , 228.5)
*       71 = U288/U240/vout (-139.5 , 287)
*       72 = U282/U238/S (-82 , 223)
*       72 = U282/Sum (-82 , 192)
*       72 = U247/CC (190.5 , 161)
*       72 = U247/U211/A (265 , 103.5)
*       74 = U282/U237/Vdd (-107.5 , 229.5)
*       74 = U282/U234/VDD (-134.5 , 228.5)
*       74 = U282/U238/VDD (-12.5 , 226)
*       75 = U279/U215/VDD (-257 , 204.5)
*       76 = U282/U237/vin (-117 , 207)
*       76 = U282/U234/OUTPUT (-128 , 215.5)
*       84 = U279/U210/C (-289.5 , 251)
*       84 = U279/U213/A (-253 , 249)
*       85 = U279/U210/A (-304 , 250.5)
*       85 = U279/AA (-304 , 256.5)
*       85 = U293/Carry (-263 , 270.5)
*       85 = U293/U238/C (-263 , 303)
*       88 = U279/U229/VDD (-446 , 255.5)
*       88 = U279/U210/VDD (-336 , 252)
*       88 = U279/U213/VDD (-217.5 , 253)
*       89 = U279/U211/VDD (-336 , 201)
*       91 = U279/U210/B (-397.5 , 248.5)
*       91 = U279/BB (-397.5 , 257)
*       91 = U279/U229/vout (-439 , 235)
*       92 = U293/Sum (-379 , 270)
*       92 = U282/U238/A (19.5 , 224.5)
*       92 = U282/AA (19.5 , 228.5)
*       92 = U293/U238/S (-379 , 301)
*       94 = U279/U228/VDD (-431.5 , 203.5)
*       95 = U309/U228/INPUTB (-450 , -62)
*       95 = U244/U228/INPUTB (-450 , -17)
*       95 = U244/Y (-448.5 , 63.5)
*       95 = U279/U228/INPUTB (-450 , 175)
*       95 = U243/U228/INPUTB (-450 , 79)
*       95 = U243/Y (-448.5 , 159.5)
*       95 = U279/Y (-448.5 , 255.5)
*       95 = U293/U234/INPUTB (-450 , 278)
*       95 = U293/Y (-448 , 307)
*       95 = Y4 (-448 , 309)
*       101 = U287/U240/vin (-706.5 , 284.5)
*       101 = U287/U239/OUT (-745 , 272.5)
*       102 = U287/U239/B (-732 , 284)
*       102 = U287/Y (-732.5 , 308)
*       102 = Y5 (-732.5 , 308)
*       102 = U310/U228/INPUTB (-734.5 , -62)
*       102 = U242/U228/INPUTB (-734.5 , -17)
*       102 = U242/Y (-733 , 63.5)
*       102 = U241/U228/INPUTB (-734.5 , 79)
*       102 = U241/Y (-733 , 159.5)
*       102 = U281/U234/INPUTB (-734.5 , 199)
*       102 = U281/Y (-732.5 , 228)
*       103 = U279/CC (-378.5 , 257)
*       103 = U279/U211/A (-304 , 199.5)
*       103 = U287/U240/vout (-721 , 286)
*       104 = U281/U237/vout (-670 , 205)
*       104 = U281/U238/B (-655.5 , 221.5)
*       106 = U299/U234/VDD (-993 , 227.5)
*       106 = U299/U232/VDD (-906.9 , 225.1)
*       106 = U281/U237/Vdd (-689 , 228.5)
*       106 = U281/U234/VDD (-716 , 227.5)
*       106 = U281/U238/VDD (-594 , 225)
*       107 = U281/U237/vin (-698.5 , 206)
*       107 = U281/U234/OUTPUT (-709.5 , 214.5)
*       115 = U299/U232/A (-874.9 , 223.6)
*       115 = U299/AA (-875 , 228.5)
*       115 = U298/Carry (-860 , 270.5)
*       115 = U298/U232/C (-860.4 , 302.1)
*       116 = U298/U234/OUTPUT (-986.5 , 292.5)
*       116 = U298/U232/B (-968.4 , 299.6)
*       117 = U299/U234/INPUTA (-1067 , 197)
*       117 = U299/X (-1072 , 211)
*       117 = X1 (-1073 , 208.5)
*       117 = U281/U234/INPUTA (-790 , 197)
*       117 = U281/X (-795 , 210.5)
*       117 = U279/U228/INPUTA (-505.5 , 173)
*       117 = U279/X (-510.5 , 212)
*       117 = U282/U234/INPUTA (-208.5 , 198)
*       117 = U282/X (-213.5 , 211.5)
*       117 = U283/U234/INPUTA (76 , 198)
*       117 = U283/X (71 , 211.5)
*       117 = U284/U234/INPUTA (360 , 198)
*       117 = U284/X (355 , 211.5)
*       117 = U285/U234/INPUTA (644.5 , 198)
*       117 = U285/X (639.5 , 211.5)
*       118 = U299/U234/OUTPUT (-986.5 , 214.5)
*       118 = U299/U232/B (-968.4 , 221.6)
*       119 = U298/Sum (-976.5 , 270)
*       119 = U281/U238/A (-562 , 223.5)
*       119 = U281/AA (-562 , 227.5)
*       119 = U298/U232/S (-976.4 , 300.1)
*       120 = U299/U232/S (-976.4 , 222.1)
*       120 = U299/Sum (-976.5 , 192)
*       120 = U241/U211/A (-588.5 , 103.5)
*       120 = U241/CC (-663 , 161)
*       122 = U251/U213/A (884.5 , 153)
*       122 = U251/U210/C (848 , 155)
*       129 = U251/U210/A (833.5 , 154.5)
*       129 = U251/AA (833.5 , 160.5)
*       129 = U285/U238/C (887 , 225)
*       129 = U285/Carry (887 , 192.5)
*       135 = U251/U229/VDD (691.5 , 159.5)
*       135 = U251/U210/VDD (801.5 , 156)
*       135 = U251/U213/VDD (920 , 157)
*       136 = U241/U228/VDD (-716 , 107.5)
*       136 = U241/U211/VDD (-620.5 , 105)
*       136 = U241/U215/VDD (-541.5 , 108.5)
*       136 = U243/U228/VDD (-431.5 , 107.5)
*       136 = U243/U211/VDD (-336 , 105)
*       136 = U243/U215/VDD (-257 , 108.5)
*       136 = U245/U228/VDD (-147 , 107.5)
*       136 = U245/U211/VDD (-51.5 , 105)
*       136 = U245/U215/VDD (27.5 , 108.5)
*       136 = U247/U228/VDD (137.5 , 107.5)
*       136 = U247/U215/VDD (312 , 108.5)
*       136 = U247/U211/VDD (233 , 105)
*       136 = U249/U228/VDD (421.5 , 107.5)
*       136 = U249/U211/VDD (517 , 105)
*       136 = U249/U215/VDD (596 , 108.5)
*       136 = U251/U228/VDD (706 , 107.5)
*       136 = U251/U211/VDD (801.5 , 105)
*       136 = U251/U215/VDD (880.5 , 108.5)
*       137 = U251/U229/vout (698.5 , 139)
*       137 = U251/U210/B (740 , 152.5)
*       137 = U251/BB (740 , 161)
*       139 = U249/U213/A (600 , 153)
*       139 = U249/U210/C (563.5 , 155)
*       151 = U249/U210/A (549 , 154.5)
*       151 = U249/AA (549 , 160.5)
*       151 = U284/U238/C (602.5 , 225)
*       151 = U284/Carry (602.5 , 192.5)
*       152 = U249/U229/vin (428.5 , 137.5)
*       152 = U249/U228/OUTPUT (428 , 94.5)
*       153 = U249/U229/vout (414 , 139)
*       153 = U249/U210/B (455.5 , 152.5)
*       153 = U249/BB (455.5 , 161)
*       156 = U249/U229/VDD (407 , 159.5)
*       156 = U249/U210/VDD (517 , 156)
*       156 = U249/U213/VDD (635.5 , 157)
*       157 = U247/U215/vin (333.5 , 86.5)
*       157 = U247/U213/O/P (345 , 145)
*       158 = U247/U213/A (316 , 153)
*       158 = U247/U210/C (279.5 , 155)
*       167 = U247/U210/B (171.5 , 152.5)
*       167 = U247/BB (171.5 , 161)
*       167 = U247/U229/vout (130 , 139)
*       168 = U247/U210/A (265 , 154.5)
*       168 = U247/AA (265 , 160.5)
*       168 = U283/U238/C (318.5 , 225)
*       168 = U283/Carry (318.5 , 192.5)
*       172 = U247/U229/vin (144.5 , 137.5)
*       172 = U247/U228/OUTPUT (144 , 94.5)
*       173 = U247/U229/VDD (123 , 159.5)
*       173 = U247/U210/VDD (233 , 156)
*       173 = U247/U213/VDD (351.5 , 157)
*       177 = U245/U210/C (-5 , 155)
*       177 = U245/U213/A (31.5 , 153)
*       178 = U245/U210/A (-19.5 , 154.5)
*       178 = U245/AA (-19.5 , 160.5)
*       178 = U282/U238/C (34 , 225)
*       178 = U282/Carry (34 , 192.5)
*       181 = U245/U229/VDD (-161.5 , 159.5)
*       181 = U245/U210/VDD (-51.5 , 156)
*       181 = U245/U213/VDD (67 , 157)
*       188 = U245/U210/B (-113 , 152.5)
*       188 = U245/BB (-113 , 161)
*       188 = U245/U229/vout (-154.5 , 139)
*       190 = U245/U229/vin (-140 , 137.5)
*       190 = U245/U228/OUTPUT (-140.5 , 94.5)
*       191 = U279/U215/vin (-235.5 , 182.5)
*       191 = U279/U213/O/P (-224 , 241)
*       200 = U279/U211/C (-289.5 , 200)
*       200 = U279/U213/B (-237.5 , 247.5)
*       201 = U243/U210/C (-289.5 , 155)
*       201 = U243/U213/A (-253 , 153)
*       202 = U243/U210/A (-304 , 154.5)
*       202 = U243/AA (-304 , 160.5)
*       202 = U279/Carry (-250.5 , 169)
*       202 = U279/U215/vout (-250 , 184)
*       207 = U243/U229/VDD (-446 , 159.5)
*       207 = U243/U210/VDD (-336 , 156)
*       207 = U243/U213/VDD (-217.5 , 157)
*       210 = U279/Sum (-405.5 , 168.5)
*       210 = U279/U211/S (-405.5 , 198)
*       210 = U245/CC (-94 , 161)
*       210 = U245/U211/A (-19.5 , 103.5)
*       211 = U243/U210/B (-397.5 , 152.5)
*       211 = U243/BB (-397.5 , 161)
*       211 = U243/U229/vout (-439 , 139)
*       213 = U279/U211/B (-397.5 , 197.5)
*       213 = U279/U210/S (-405.5 , 249)
*       214 = U279/U229/vin (-424.5 , 233.5)
*       214 = U279/U228/OUTPUT (-425 , 190.5)
*       215 = U243/U229/vin (-424.5 , 137.5)
*       215 = U243/U228/OUTPUT (-425 , 94.5)
*       225 = U241/U210/C (-574 , 155)
*       225 = U241/U213/A (-537.5 , 153)
*       226 = U243/CC (-378.5 , 161)
*       226 = U243/U211/A (-304 , 103.5)
*       226 = U281/U238/S (-663.5 , 222)
*       226 = U281/Sum (-663.5 , 191)
*       227 = U241/U210/A (-588.5 , 154.5)
*       227 = U241/AA (-588.5 , 160.5)
*       227 = U281/U238/C (-547.5 , 224)
*       227 = U281/Carry (-547.5 , 191.5)
*       228 = U241/U229/VDD (-730.5 , 159.5)
*       228 = U241/U210/VDD (-620.5 , 156)
*       228 = U241/U213/VDD (-502 , 157)
*       231 = U241/U210/B (-682 , 152.5)
*       231 = U241/BB (-682 , 161)
*       231 = U241/U229/vout (-723.5 , 139)
*       233 = U241/U229/vin (-709 , 137.5)
*       233 = U241/U228/OUTPUT (-709.5 , 94.5)
*       239 = U300/U232/A (-874.9 , 128.6)
*       239 = U300/AA (-875 , 133.5)
*       239 = U299/U232/C (-860.4 , 224.1)
*       239 = U299/Carry (-860 , 192.5)
*       240 = U300/U234/VDD (-993 , 132.5)
*       240 = U300/U232/VDD (-906.9 , 130.1)
*       241 = U300/U234/INPUTA (-1067 , 102)
*       241 = U300/X (-1072 , 116)
*       241 = X2 (-1073 , 113.5)
*       241 = U241/U228/INPUTA (-790 , 77)
*       241 = U241/X (-795 , 116)
*       241 = U243/U228/INPUTA (-505.5 , 77)
*       241 = U243/X (-510.5 , 116)
*       241 = U245/U228/INPUTA (-221 , 77)
*       241 = U245/X (-226 , 116)
*       241 = U247/U228/INPUTA (63.5 , 77)
*       241 = U247/X (58.5 , 116)
*       241 = U249/U228/INPUTA (347.5 , 77)
*       241 = U249/X (342.5 , 116)
*       241 = U251/U228/INPUTA (632 , 77)
*       241 = U251/X (627 , 116)
*       242 = U300/U234/OUTPUT (-986.5 , 119.5)
*       242 = U300/U232/B (-968.4 , 126.6)
*       243 = U300/U232/S (-976.4 , 127.1)
*       243 = U300/Sum (-976.5 , 97)
*       243 = U242/U211/A (-588.5 , 7.5)
*       243 = U242/CC (-663 , 65)
*       245 = U251/U215/vin (902 , 86.5)
*       245 = U251/U213/O/P (913.5 , 145)
*       246 = U252/U213/A (884.5 , 57)
*       246 = U252/U210/C (848 , 59)
*       247 = U251/U213/B (900 , 151.5)
*       247 = U251/U211/C (848 , 104)
*       254 = U252/U210/A (833.5 , 58.5)
*       254 = U252/AA (833.5 , 64.5)
*       254 = U251/Carry (887 , 73)
*       254 = U251/U215/vout (887.5 , 88)
*       260 = U251/U211/B (740 , 101.5)
*       260 = U251/U210/S (732 , 153)
*       261 = U251/Sum (732 , 72.5)
*       261 = U251/U211/S (732 , 102)
*       261 = P2 (922 , 99.5)
*       262 = U251/U229/vin (713 , 137.5)
*       262 = U251/U228/OUTPUT (712.5 , 94.5)
*       263 = U242/U228/VDD (-716 , 11.5)
*       263 = U242/U211/VDD (-620.5 , 9)
*       263 = U242/U215/VDD (-541.5 , 12.5)
*       263 = U244/U228/VDD (-431.5 , 11.5)
*       263 = U244/U211/VDD (-336 , 9)
*       263 = U244/U215/VDD (-257 , 12.5)
*       263 = U246/U228/VDD (-147 , 11.5)
*       263 = U246/U211/VDD (-51.5 , 9)
*       263 = U246/U215/VDD (27.5 , 12.5)
*       263 = U248/U228/VDD (137.5 , 11.5)
*       263 = U248/U215/VDD (312 , 12.5)
*       263 = U248/U211/VDD (233 , 9)
*       263 = U250/U228/VDD (421.5 , 11.5)
*       263 = U250/U211/VDD (517 , 9)
*       263 = U250/U215/VDD (596 , 12.5)
*       263 = U252/U228/VDD (706 , 11.5)
*       263 = U252/U211/VDD (801.5 , 9)
*       263 = U252/U215/VDD (880.5 , 12.5)
*       264 = U252/U229/vout (698.5 , 43)
*       264 = U252/U210/B (740 , 56.5)
*       264 = U252/BB (740 , 65)
*       266 = U249/U215/vin (617.5 , 86.5)
*       266 = U249/U213/O/P (629 , 145)
*       267 = U250/U213/A (600 , 57)
*       267 = U250/U210/C (563.5 , 59)
*       268 = U249/U213/B (615.5 , 151.5)
*       268 = U249/U211/C (563.5 , 104)
*       280 = U249/U211/B (455.5 , 101.5)
*       280 = U249/U210/S (447.5 , 153)
*       281 = U249/Sum (447.5 , 72.5)
*       281 = U249/U211/S (447.5 , 102)
*       281 = U252/CC (759 , 65)
*       281 = U252/U211/A (833.5 , 7.5)
*       282 = U250/U210/A (549 , 58.5)
*       282 = U250/AA (549 , 64.5)
*       282 = U249/Carry (602.5 , 73)
*       282 = U249/U215/vout (603 , 88)
*       283 = U250/U229/vin (428.5 , 41.5)
*       283 = U250/U228/OUTPUT (428 , -1.5)
*       284 = U250/U229/vout (414 , 43)
*       284 = U250/U210/B (455.5 , 56.5)
*       284 = U250/BB (455.5 , 65)
*       287 = U242/U229/VDD (-730.5 , 63.5)
*       287 = U242/U210/VDD (-620.5 , 60)
*       287 = U242/U213/VDD (-502 , 61)
*       287 = U244/U229/VDD (-446 , 63.5)
*       287 = U244/U210/VDD (-336 , 60)
*       287 = U244/U213/VDD (-217.5 , 61)
*       287 = U246/U229/VDD (-161.5 , 63.5)
*       287 = U246/U210/VDD (-51.5 , 60)
*       287 = U248/U229/VDD (123 , 63.5)
*       287 = U246/U213/VDD (67 , 61)
*       287 = U248/U210/VDD (233 , 60)
*       287 = U250/U229/VDD (407 , 63.5)
*       287 = U248/U213/VDD (351.5 , 61)
*       287 = U250/U210/VDD (517 , 60)
*       287 = U252/U229/VDD (691.5 , 63.5)
*       287 = U250/U213/VDD (635.5 , 61)
*       287 = U252/U210/VDD (801.5 , 60)
*       287 = U252/U213/VDD (920 , 61)
*       288 = U248/U215/vin (333.5 , -9.5)
*       288 = U248/U213/O/P (345 , 49)
*       289 = U248/U213/A (316 , 57)
*       289 = U248/U210/C (279.5 , 59)
*       290 = U247/U211/C (279.5 , 104)
*       290 = U247/U213/B (331.5 , 151.5)
*       299 = U247/U211/B (171.5 , 101.5)
*       299 = U247/U210/S (163.5 , 153)
*       300 = U247/Sum (163.5 , 72.5)
*       300 = U247/U211/S (163.5 , 102)
*       300 = U250/CC (474.5 , 65)
*       300 = U250/U211/A (549 , 7.5)
*       301 = U248/U210/B (171.5 , 56.5)
*       301 = U248/BB (171.5 , 65)
*       301 = U248/U229/vout (130 , 43)
*       302 = U248/U210/A (265 , 58.5)
*       302 = U248/AA (265 , 64.5)
*       302 = U247/Carry (318.5 , 73)
*       302 = U247/U215/vout (319 , 88)
*       306 = U245/U215/vin (49 , 86.5)
*       306 = U245/U213/O/P (60.5 , 145)
*       307 = U248/U229/vin (144.5 , 41.5)
*       307 = U248/U228/OUTPUT (144 , -1.5)
*       311 = U246/U210/C (-5 , 59)
*       311 = U246/U213/A (31.5 , 57)
*       312 = U245/U211/C (-5 , 104)
*       312 = U245/U213/B (47 , 151.5)
*       313 = U246/U210/A (-19.5 , 58.5)
*       313 = U246/AA (-19.5 , 64.5)
*       313 = U245/Carry (34 , 73)
*       313 = U245/U215/vout (34.5 , 88)
*       322 = U245/U211/B (-113 , 101.5)
*       322 = U245/U210/S (-121 , 153)
*       323 = U245/Sum (-121 , 72.5)
*       323 = U245/U211/S (-121 , 102)
*       323 = U248/CC (190.5 , 65)
*       323 = U248/U211/A (265 , 7.5)
*       324 = U246/U210/B (-113 , 56.5)
*       324 = U246/BB (-113 , 65)
*       324 = U246/U229/vout (-154.5 , 43)
*       326 = U243/U215/vin (-235.5 , 86.5)
*       326 = U243/U213/O/P (-224 , 145)
*       327 = U246/U229/vin (-140 , 41.5)
*       327 = U246/U228/OUTPUT (-140.5 , -1.5)
*       335 = U244/U210/C (-289.5 , 59)
*       335 = U244/U213/A (-253 , 57)
*       336 = U243/U211/C (-289.5 , 104)
*       336 = U243/U213/B (-237.5 , 151.5)
*       337 = U244/U210/A (-304 , 58.5)
*       337 = U244/AA (-304 , 64.5)
*       337 = U243/Carry (-250.5 , 73)
*       337 = U243/U215/vout (-250 , 88)
*       342 = U243/U211/B (-397.5 , 101.5)
*       342 = U243/U210/S (-405.5 , 153)
*       343 = U243/Sum (-405.5 , 72.5)
*       343 = U243/U211/S (-405.5 , 102)
*       343 = U246/CC (-94 , 65)
*       343 = U246/U211/A (-19.5 , 7.5)
*       344 = U244/U210/B (-397.5 , 56.5)
*       344 = U244/BB (-397.5 , 65)
*       344 = U244/U229/vout (-439 , 43)
*       346 = U241/U215/vin (-520 , 86.5)
*       346 = U241/U213/O/P (-508.5 , 145)
*       347 = U244/U229/vin (-424.5 , 41.5)
*       347 = U244/U228/OUTPUT (-425 , -1.5)
*       357 = U242/U210/C (-574 , 59)
*       357 = U242/U213/A (-537.5 , 57)
*       358 = U241/U211/C (-574 , 104)
*       358 = U241/U213/B (-522 , 151.5)
*       359 = U242/U210/A (-588.5 , 58.5)
*       359 = U242/AA (-588.5 , 64.5)
*       359 = U241/Carry (-535 , 73)
*       359 = U241/U215/vout (-534.5 , 88)
*       362 = U241/U211/B (-682 , 101.5)
*       362 = U241/U210/S (-690 , 153)
*       363 = U241/Sum (-690 , 72.5)
*       363 = U241/U211/S (-690 , 102)
*       363 = U244/CC (-378.5 , 65)
*       363 = U244/U211/A (-304 , 7.5)
*       364 = U242/U210/B (-682 , 56.5)
*       364 = U242/BB (-682 , 65)
*       364 = U242/U229/vout (-723.5 , 43)
*       366 = U242/U229/vin (-709 , 41.5)
*       366 = U242/U228/OUTPUT (-709.5 , -1.5)
*       372 = U301/U232/A (-874.9 , 32.6)
*       372 = U301/AA (-875 , 37.5)
*       372 = U300/U232/C (-860.4 , 129.1)
*       372 = U300/Carry (-860 , 97.5)
*       373 = U301/U234/VDD (-993 , 36.5)
*       373 = U301/U232/VDD (-906.9 , 34.1)
*       374 = U301/U234/INPUTA (-1067 , 6)
*       374 = U301/X (-1072 , 20)
*       374 = X3 (-1073 , 17.5)
*       374 = U242/U228/INPUTA (-790 , -19)
*       374 = U242/X (-795 , 20)
*       374 = U244/U228/INPUTA (-505.5 , -19)
*       374 = U244/X (-510.5 , 20)
*       374 = U246/U228/INPUTA (-221 , -19)
*       374 = U246/X (-226 , 20)
*       374 = U248/U228/INPUTA (63.5 , -19)
*       374 = U248/X (58.5 , 20)
*       374 = U250/U228/INPUTA (347.5 , -19)
*       374 = U250/X (342.5 , 20)
*       374 = U252/U228/INPUTA (632 , -19)
*       374 = U252/X (627 , 20)
*       375 = U301/U234/OUTPUT (-986.5 , 23.5)
*       375 = U301/U232/B (-968.4 , 30.6)
*       376 = U301/U232/S (-976.4 , 31.1)
*       376 = U301/Sum (-976.5 , 1)
*       376 = U310/U211/A (-598 , -88.5)
*       376 = U310/CC (-672.5 , -31)
*       378 = U294/U215/vin (892.5 , -105.5)
*       378 = U294/U213/O/P (904 , -47)
*       379 = U294/U213/A (875 , -39)
*       379 = U294/U210/C (838.5 , -37)
*       380 = U294/U213/B (890.5 , -40.5)
*       380 = U294/U211/C (838.5 , -88)
*       381 = U252/U215/vin (902 , -9.5)
*       381 = U252/U213/O/P (913.5 , 49)
*       382 = U252/U213/B (900 , 55.5)
*       382 = U252/U211/C (848 , 8)
*       394 = U252/U211/B (740 , 5.5)
*       394 = U252/U210/S (732 , 57)
*       395 = U252/U211/S (732 , 6)
*       395 = U252/Sum (732 , -23.5)
*       395 = P3 (922 , 3.5)
*       396 = U294/U210/A (824 , -37.5)
*       396 = U294/AA (824 , -31.5)
*       396 = U252/U215/vout (887.5 , -8)
*       396 = U252/Carry (887 , -23)
*       397 = U294/U210/S (722.5 , -39)
*       397 = U294/U211/B (730.5 , -90.5)
*       398 = U252/U229/vin (713 , 41.5)
*       398 = U252/U228/OUTPUT (712.5 , -1.5)
*       399 = U310/U211/VDD (-630 , -87)
*       399 = U310/U215/VDD (-551 , -83.5)
*       399 = U309/U211/VDD (-345.5 , -87)
*       399 = U309/U215/VDD (-266.5 , -83.5)
*       399 = U308/U215/VDD (18 , -83.5)
*       399 = U308/U211/VDD (-61 , -87)
*       399 = U297/U211/VDD (223.5 , -87)
*       399 = U297/U215/VDD (302.5 , -83.5)
*       399 = U295/U211/VDD (507.5 , -87)
*       399 = U295/U215/VDD (586.5 , -83.5)
*       399 = U294/U211/VDD (792 , -87)
*       399 = U294/U215/VDD (871 , -83.5)
*       400 = U310/U228/VDD (-716 , -33.5)
*       400 = U310/U210/VDD (-630 , -36)
*       400 = U310/U213/VDD (-511.5 , -35)
*       400 = U309/U228/VDD (-431.5 , -33.5)
*       400 = U309/U210/VDD (-345.5 , -36)
*       400 = U309/U213/VDD (-227 , -35)
*       400 = U308/U228/VDD (-147 , -33.5)
*       400 = U308/U210/VDD (-61 , -36)
*       400 = U308/U213/VDD (57.5 , -35)
*       400 = U297/U228/VDD (137.5 , -33.5)
*       400 = U297/U210/VDD (223.5 , -36)
*       400 = U297/U213/VDD (342 , -35)
*       400 = U295/U228/VDD (421.5 , -33.5)
*       400 = U295/U210/VDD (507.5 , -36)
*       400 = U295/U213/VDD (626 , -35)
*       400 = U294/U228/VDD (706 , -33.5)
*       400 = U294/U210/VDD (792 , -36)
*       400 = U294/U213/VDD (910.5 , -35)
*       401 = U294/U228/OUTPUT (712.5 , -46.5)
*       401 = U294/U210/B (730.5 , -39.5)
*       401 = U294/BB (730.5 , -31)
*       402 = U294/U211/S (722.5 , -90)
*       402 = U294/Sum (722.5 , -119.5)
*       402 = P4 (912.5 , -92.5)
*       404 = U295/U215/vin (608 , -105.5)
*       404 = U295/U213/O/P (619.5 , -47)
*       405 = U295/U213/A (590.5 , -39)
*       405 = U295/U210/C (554 , -37)
*       406 = U295/U213/B (606 , -40.5)
*       406 = U295/U211/C (554 , -88)
*       407 = U250/U215/vin (617.5 , -9.5)
*       407 = U250/U213/O/P (629 , 49)
*       408 = U250/U213/B (615.5 , 55.5)
*       408 = U250/U211/C (563.5 , 8)
*       419 = U295/U211/B (446 , -90.5)
*       419 = U295/U210/S (438 , -39)
*       421 = U250/U211/B (455.5 , 5.5)
*       421 = U250/U210/S (447.5 , 57)
*       422 = U250/U211/S (447.5 , 6)
*       422 = U250/Sum (447.5 , -23.5)
*       422 = U294/U211/A (824 , -88.5)
*       422 = U294/CC (749.5 , -31)
*       423 = U295/U211/S (438 , -90)
*       423 = U295/Sum (438 , -119.5)
*       423 = U269/B (730.5 , -141.5)
*       424 = U295/U210/A (539.5 , -37.5)
*       424 = U295/AA (539.5 , -31.5)
*       424 = U250/U215/vout (603 , -8)
*       424 = U250/Carry (602.5 , -23)
*       425 = U295/U210/B (446 , -39.5)
*       425 = U295/BB (446 , -31)
*       425 = U295/U228/OUTPUT (428 , -46.5)
*       427 = U297/U215/vin (324 , -105.5)
*       427 = U297/U213/O/P (335.5 , -47)
*       428 = U297/U213/A (306.5 , -39)
*       428 = U297/U210/C (270 , -37)
*       429 = U297/U213/B (322 , -40.5)
*       429 = U297/U211/C (270 , -88)
*       430 = U248/U211/C (279.5 , 8)
*       430 = U248/U213/B (331.5 , 55.5)
*       441 = U297/U211/B (162 , -90.5)
*       441 = U297/U210/S (154 , -39)
*       443 = U248/U211/B (171.5 , 5.5)
*       443 = U248/U210/S (163.5 , 57)
*       444 = U248/U211/S (163.5 , 6)
*       444 = U248/Sum (163.5 , -23.5)
*       444 = U295/CC (465 , -31)
*       444 = U295/U211/A (539.5 , -88.5)
*       445 = U297/U211/S (154 , -90)
*       445 = U297/Sum (154 , -119.5)
*       445 = U296/U210/B (446 , -141.5)
*       445 = U296/BB (446 , -133)
*       446 = U297/U210/A (255.5 , -37.5)
*       446 = U297/AA (255.5 , -31.5)
*       446 = U248/U215/vout (319 , -8)
*       446 = U248/Carry (318.5 , -23)
*       448 = U308/U215/vin (39.5 , -105.5)
*       448 = U308/U213/O/P (51 , -47)
*       449 = U297/U210/B (162 , -39.5)
*       449 = U297/BB (162 , -31)
*       449 = U297/U228/OUTPUT (144 , -46.5)
*       450 = U246/U215/vin (49 , -9.5)
*       450 = U246/U213/O/P (60.5 , 49)
*       452 = U308/U213/A (22 , -39)
*       452 = U308/U210/C (-14.5 , -37)
*       453 = U308/U211/C (-14.5 , -88)
*       453 = U308/U213/B (37.5 , -40.5)
*       454 = U246/U211/C (-5 , 8)
*       454 = U246/U213/B (47 , 55.5)
*       458 = U308/U211/B (-122.5 , -90.5)
*       458 = U308/U210/S (-130.5 , -39)
*       460 = U246/U211/B (-113 , 5.5)
*       460 = U246/U210/S (-121 , 57)
*       461 = U246/U211/S (-121 , 6)
*       461 = U246/Sum (-121 , -23.5)
*       461 = U297/CC (181 , -31)
*       461 = U297/U211/A (255.5 , -88.5)
*       462 = U308/U211/S (-130.5 , -90)
*       462 = U308/Sum (-130.5 , -119.5)
*       462 = U307/U210/B (162 , -141.5)
*       462 = U307/BB (162 , -133)
*       464 = U308/U210/A (-29 , -37.5)
*       464 = U308/AA (-29 , -31.5)
*       464 = U246/U215/vout (34.5 , -8)
*       464 = U246/Carry (34 , -23)
*       471 = U309/U215/vin (-245 , -105.5)
*       471 = U309/U213/O/P (-233.5 , -47)
*       472 = U308/U210/B (-122.5 , -39.5)
*       472 = U308/BB (-122.5 , -31)
*       472 = U308/U228/OUTPUT (-140.5 , -46.5)
*       473 = U244/U215/vin (-235.5 , -9.5)
*       473 = U244/U213/O/P (-224 , 49)
*       477 = U309/U211/C (-299 , -88)
*       477 = U309/U213/B (-247 , -40.5)
*       478 = U309/U210/C (-299 , -37)
*       478 = U309/U213/A (-262.5 , -39)
*       479 = U244/U211/C (-289.5 , 8)
*       479 = U244/U213/B (-237.5 , 55.5)
*       480 = U309/U210/A (-313.5 , -37.5)
*       480 = U309/AA (-313.5 , -31.5)
*       480 = U244/U215/vout (-250 , -8)
*       480 = U244/Carry (-250.5 , -23)
*       487 = U309/U211/B (-407 , -90.5)
*       487 = U309/U210/S (-415 , -39)
*       488 = U244/U211/B (-397.5 , 5.5)
*       488 = U244/U210/S (-405.5 , 57)
*       489 = U244/U211/S (-405.5 , 6)
*       489 = U244/Sum (-405.5 , -23.5)
*       489 = U308/CC (-103.5 , -31)
*       489 = U308/U211/A (-29 , -88.5)
*       490 = U309/U211/S (-415 , -90)
*       490 = U309/Sum (-415 , -119.5)
*       490 = U306/U210/B (-122.5 , -141.5)
*       490 = U306/BB (-122.5 , -133)
*       494 = U310/U215/vin (-529.5 , -105.5)
*       494 = U310/U213/O/P (-518 , -47)
*       495 = U309/U210/B (-407 , -39.5)
*       495 = U309/BB (-407 , -31)
*       495 = U309/U228/OUTPUT (-425 , -46.5)
*       496 = U242/U215/vin (-520 , -9.5)
*       496 = U242/U213/O/P (-508.5 , 49)
*       504 = U310/U211/C (-583.5 , -88)
*       504 = U310/U213/B (-531.5 , -40.5)
*       505 = U310/U210/C (-583.5 , -37)
*       505 = U310/U213/A (-547 , -39)
*       506 = U242/U211/C (-574 , 8)
*       506 = U242/U213/B (-522 , 55.5)
*       507 = U310/U210/A (-598 , -37.5)
*       507 = U310/AA (-598 , -31.5)
*       507 = U242/U215/vout (-534.5 , -8)
*       507 = U242/Carry (-535 , -23)
*       512 = U310/U211/B (-691.5 , -90.5)
*       512 = U310/U210/S (-699.5 , -39)
*       513 = U242/U211/B (-682 , 5.5)
*       513 = U242/U210/S (-690 , 57)
*       514 = U242/U211/S (-690 , 6)
*       514 = U242/Sum (-690 , -23.5)
*       514 = U309/CC (-388 , -31)
*       514 = U309/U211/A (-313.5 , -88.5)
*       515 = U310/U211/S (-699.5 , -90)
*       515 = U310/Sum (-699.5 , -119.5)
*       515 = U305/U210/B (-407 , -141.5)
*       515 = U305/BB (-407 , -133)
*       518 = U310/U210/B (-691.5 , -39.5)
*       518 = U310/BB (-691.5 , -31)
*       518 = U310/U228/OUTPUT (-709.5 , -46.5)
*       522 = U302/U237/vout (-947 , -81)
*       522 = U302/U238/B (-932.5 , -64.5)
*       523 = U302/U238/S (-940.5 , -64)
*       523 = U302/Sum (-940.5 , -95)
*       523 = U304/U210/B (-691.5 , -141.5)
*       523 = U304/BB (-691.5 , -133)
*       524 = U302/U238/A (-839 , -62.5)
*       524 = U302/AA (-839 , -58.5)
*       524 = U301/U232/C (-860.4 , 33.1)
*       524 = U301/Carry (-860 , 1.5)
*       526 = U302/U234/INPUTB (-1011.5 , -87)
*       526 = U302/Y (-1009.5 , -58)
*       526 = U301/U234/INPUTB (-1011.5 , 8)
*       526 = U301/Y (-1009.5 , 37)
*       526 = U300/U234/INPUTB (-1011.5 , 104)
*       526 = U300/Y (-1009.5 , 133)
*       526 = U299/U234/INPUTB (-1011.5 , 199)
*       526 = U299/Y (-1009.5 , 228)
*       526 = U298/U234/INPUTB (-1011.5 , 277)
*       526 = U298/Y (-1009.5 , 306)
*       526 = Y6 (-1009.5 , 308)
*       527 = U302/U237/Vdd (-966 , -57.5)
*       527 = U302/U234/VDD (-993 , -58.5)
*       527 = U302/U238/VDD (-871 , -61)
*       528 = U302/U234/INPUTA (-1067 , -89)
*       528 = U302/X (-1072 , -75.5)
*       528 = X4 (-1073 , -77.5)
*       528 = U310/U228/INPUTA (-790 , -64)
*       528 = U310/X (-795 , -76)
*       528 = U309/U228/INPUTA (-505.5 , -64)
*       528 = U309/X (-510.5 , -76)
*       528 = U308/U228/INPUTA (-221 , -64)
*       528 = U308/X (-226 , -76)
*       528 = U297/U228/INPUTA (63.5 , -64)
*       528 = U297/X (58.5 , -76)
*       528 = U295/U228/INPUTA (347.5 , -64)
*       528 = U295/X (342.5 , -76)
*       528 = U294/U228/INPUTA (632 , -64)
*       528 = U294/X (627 , -76)
*       529 = U302/U237/vin (-975.5 , -80)
*       529 = U302/U234/OUTPUT (-986.5 , -71.5)
*       536 = U269/A (824 , -139.5)
*       536 = U294/U215/vout (878 , -104)
*       536 = U294/Carry (877.5 , -119)
*       537 = U303/U210/B (-989 , -141.5)
*       537 = U303/BB (-989 , -133)
*       537 = U303/U210/VDD (-927.5 , -138)
*       537 = U303/U213/VDD (-809 , -137)
*       537 = U304/U210/VDD (-630 , -138)
*       537 = U304/U213/VDD (-511.5 , -137)
*       537 = U305/U210/VDD (-345.5 , -138)
*       537 = U305/U213/VDD (-227 , -137)
*       537 = U306/U210/VDD (-61 , -138)
*       537 = U306/U213/VDD (57.5 , -137)
*       537 = U307/U210/VDD (223.5 , -138)
*       537 = U307/U213/VDD (342 , -137)
*       537 = U296/U210/VDD (507.5 , -138)
*       537 = U296/U213/VDD (626 , -137)
*       537 = U269/VDD (792 , -138)
*       538 = U269/S (722.5 , -141)
*       538 = P5 (912.5 , -145.5)
*       539 = U296/U215/vin (608 , -207.5)
*       539 = U296/U213/O/P (619.5 , -149)
*       540 = U296/U213/A (590.5 , -141)
*       540 = U296/U210/C (554 , -139)
*       541 = U296/U213/B (606 , -142.5)
*       541 = U296/U211/C (554 , -190)
*       552 = U296/U211/B (446 , -192.5)
*       552 = U296/U210/S (438 , -141)
*       553 = U296/U211/S (438 , -192)
*       553 = U296/Sum (438 , -221.5)
*       553 = P6 (438 , -223)
*       555 = U296/CC (465 , -133)
*       555 = U296/U211/A (539.5 , -190.5)
*       555 = U269/C (838.5 , -139)
*       556 = U296/U210/A (539.5 , -139.5)
*       556 = U296/AA (539.5 , -133.5)
*       556 = U295/U215/vout (593.5 , -104)
*       556 = U295/Carry (593 , -119)
*       557 = U303/U215/VDD (-848.5 , -185.5)
*       557 = U304/U211/VDD (-630 , -189)
*       557 = U304/U215/VDD (-551 , -185.5)
*       557 = U305/U211/VDD (-345.5 , -189)
*       557 = U305/U215/VDD (-266.5 , -185.5)
*       557 = U306/U215/VDD (18 , -185.5)
*       557 = U306/U211/VDD (-61 , -189)
*       557 = U307/U211/VDD (223.5 , -189)
*       557 = U307/U215/VDD (302.5 , -185.5)
*       557 = U296/U211/VDD (507.5 , -189)
*       557 = U296/U215/VDD (586.5 , -185.5)
*       558 = U307/U215/vin (324 , -207.5)
*       558 = U307/U213/O/P (335.5 , -149)
*       559 = U307/U213/A (306.5 , -141)
*       559 = U307/U210/C (270 , -139)
*       560 = U307/U213/B (322 , -142.5)
*       560 = U307/U211/C (270 , -190)
*       571 = U307/U211/B (162 , -192.5)
*       571 = U307/U210/S (154 , -141)
*       572 = U307/U211/S (154 , -192)
*       572 = U307/Sum (154 , -221.5)
*       572 = P7 (154 , -223)
*       574 = U307/U210/A (255.5 , -139.5)
*       574 = U307/AA (255.5 , -133.5)
*       574 = U297/U215/vout (309.5 , -104)
*       574 = U297/Carry (309 , -119)
*       575 = U307/CC (181 , -133)
*       575 = U307/U211/A (255.5 , -190.5)
*       575 = U296/U215/vout (593.5 , -206)
*       575 = U296/Carry (593 , -221)
*       576 = U306/U215/vin (39.5 , -207.5)
*       576 = U306/U213/O/P (51 , -149)
*       578 = U306/U213/A (22 , -141)
*       578 = U306/U210/C (-14.5 , -139)
*       579 = U306/U211/C (-14.5 , -190)
*       579 = U306/U213/B (37.5 , -142.5)
*       583 = U306/U211/B (-122.5 , -192.5)
*       583 = U306/U210/S (-130.5 , -141)
*       584 = U306/U211/S (-130.5 , -192)
*       584 = U306/Sum (-130.5 , -221.5)
*       584 = P8 (-130.5 , -223)
*       587 = U306/U210/A (-29 , -139.5)
*       587 = U306/AA (-29 , -133.5)
*       587 = U308/U215/vout (25 , -104)
*       587 = U308/Carry (24.5 , -119)
*       589 = U306/CC (-103.5 , -133)
*       589 = U306/U211/A (-29 , -190.5)
*       589 = U307/U215/vout (309.5 , -206)
*       589 = U307/Carry (309 , -221)
*       594 = U305/U215/vin (-245 , -207.5)
*       594 = U305/U213/O/P (-233.5 , -149)
*       598 = U305/U211/C (-299 , -190)
*       598 = U305/U213/B (-247 , -142.5)
*       599 = U305/U210/C (-299 , -139)
*       599 = U305/U213/A (-262.5 , -141)
*       600 = U305/U210/A (-313.5 , -139.5)
*       600 = U305/AA (-313.5 , -133.5)
*       600 = U309/U215/vout (-259.5 , -104)
*       600 = U309/Carry (-260 , -119)
*       607 = U305/U211/B (-407 , -192.5)
*       607 = U305/U210/S (-415 , -141)
*       608 = U305/U211/S (-415 , -192)
*       608 = U305/Sum (-415 , -221.5)
*       608 = P9 (-415 , -223)
*       609 = U305/CC (-388 , -133)
*       609 = U305/U211/A (-313.5 , -190.5)
*       609 = U306/U215/vout (25 , -206)
*       609 = U306/Carry (24.5 , -221)
*       612 = U304/U215/vin (-529.5 , -207.5)
*       612 = U304/U213/O/P (-518 , -149)
*       620 = U304/U211/C (-583.5 , -190)
*       620 = U304/U213/B (-531.5 , -142.5)
*       621 = U304/U210/C (-583.5 , -139)
*       621 = U304/U213/A (-547 , -141)
*       622 = U304/U210/A (-598 , -139.5)
*       622 = U304/AA (-598 , -133.5)
*       622 = U310/U215/vout (-544 , -104)
*       622 = U310/Carry (-544.5 , -119)
*       627 = U304/U211/B (-691.5 , -192.5)
*       627 = U304/U210/S (-699.5 , -141)
*       628 = U304/U211/S (-699.5 , -192)
*       628 = U304/Sum (-699.5 , -221.5)
*       628 = P10 (-699.5 , -223)
*       629 = U304/U211/A (-598 , -190.5)
*       629 = U304/CC (-672.5 , -133)
*       629 = U305/U215/vout (-259.5 , -206)
*       629 = U305/Carry (-260 , -221)
*       630 = U303/U215/vin (-827 , -207.5)
*       630 = U303/U213/O/P (-815.5 , -149)
*       631 = U303/U215/vout (-841.5 , -206)
*       631 = U303/Carry (-842 , -221)
*       639 = U303/U211/C (-881 , -190)
*       639 = U303/U213/B (-829 , -142.5)
*       640 = U303/U211/A (-895.5 , -190.5)
*       640 = U303/CC (-970 , -133)
*       640 = U302/U238/C (-824.5 , -62)
*       640 = U302/Carry (-824.5 , -94.5)
*       641 = U303/U210/C (-881 , -139)
*       641 = U303/U213/A (-844.5 , -141)
*       642 = U303/U210/A (-895.5 , -139.5)
*       642 = U303/AA (-895.5 , -133.5)
*       642 = U304/U215/vout (-544 , -206)
*       642 = U304/Carry (-544.5 , -221)
*       647 = U303/U211/B (-989 , -192.5)
*       647 = U303/U210/S (-997 , -141)
*       648 = U303/U211/S (-997 , -192)
*       648 = U303/Sum (-997 , -221.5)
*       648 = P11 (-997 , -223)
*       649 = U303/U211/VDD (-927.5 , -189)



M1425 1 34 36 1 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1424 1 33 34 1 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1423 34 9 1 1 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1422 31 34 36 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1421 34 33 2 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1420 2 9 31 31 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1419 are shorted:
* D1419 1 1 D_lateral AREA=3.125E-016    $ (701.5 296.5 701.501 301.5)CMOSN1419 1 1 D_lateral AREA=3.125E-016    
M1418 3 47 4 3 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1417 31 47 4 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1416 3 46 47 3 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1415 47 9 3 3 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1414 47 46 5 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1413 5 9 31 31 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1412 are shorted:
* D1412 3 3 D_lateral AREA=3.125E-016    $ (417 296.5 417.001 301.5)CMOSN1412 3 3 D_lateral AREA=3.125E-016    
M1411 7 61 56 7 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1409 31 61 56 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
* Pins of element D1408 are shorted:
* D1408 7 7 D_lateral AREA=3.125E-016    $ (133 296.5 133.001 301.5)CMOSN1408 7 7 D_lateral AREA=3.125E-016    
M1407 61 60 7 7 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1406 61 9 7 7 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1405 61 60 6 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1404 6 9 31 31 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1403 10 68 71 10 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1402 10 69 68 10 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1401 68 9 10 10 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1400 31 68 71 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1399 68 69 8 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1398 31 9 8 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
* Pins of element D1397 are shorted:
* D1397 10 10 D_lateral AREA=3.125E-016    $ (-151.5 296.5 -151.499 301.5)CMOSN1397 10 10 D_lateral AREA=3.125E-016    
M1396 11 83 85 16 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1395 16 82 11 16 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1394 85 83 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1393 31 82 85 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1392 83 16 16 16 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1391 16 16 13 16 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1390 13 14 16 16 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1389 16 14 82 16 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1388 13 82 92 16 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1387 13 83 92 16 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1386 83 16 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1385 12 14 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1384 31 14 82 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1383 92 82 12 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1382 31 83 12 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1381 12 16 92 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1380 14 17 16 16 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1379 14 17 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1378 15 9 17 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1377 31 95 15 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1376 16 95 17 16 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1375 17 9 16 16 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1374 22 101 103 22 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1373 22 102 101 22 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1372 101 9 22 22 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1371 31 101 103 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1370 101 102 18 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1369 18 9 31 31 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
* Pins of element D1368 are shorted:
* D1368 22 22 D_lateral AREA=3.125E-016    $ (-733 295.5 -732.999 300.5)CMOSN1368 22 22 D_lateral AREA=3.125E-016    
M1367 19 112 115 22 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1366 22 113 19 22 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1365 115 112 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1364 31 113 115 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1363 112 22 22 22 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1362 22 22 21 22 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1361 21 116 22 22 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1360 22 116 113 22 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1359 21 113 119 22 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1358 21 112 119 22 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1357 112 22 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1356 31 116 20 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M1355 31 116 113 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1354 119 113 20 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1353 31 112 20 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1352 20 22 119 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1351 22 526 116 22 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1350 116 9 22 22 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1349 23 9 116 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1348 31 526 23 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1347 32 27 24 32 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1346 24 30 129 32 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1345 30 4 32 32 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1344 32 4 26 32 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1342 31 27 129 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1341 129 30 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1340 30 4 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1338 31 30 25 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1337 26 28 32 32 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1336 32 28 27 32 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1335 26 27 29 32 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1334 29 30 26 32 CMOSP L=750n W=750n AD=7.4375p PD=19.125u AS=1.109375p PS=3.375u    
M1333 28 35 32 32 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1332 25 28 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1331 31 28 27 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1330 25 27 29 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1329 29 4 25 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=1.15625p PS=3.5u    
M1328 28 35 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1327 32 33 35 32 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1326 35 117 32 32 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1325 37 117 35 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1324 31 33 37 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1323 are shorted:
* D1323 31 31 D_lateral AREA=3.125E-016    $ (709 198 714 198.001)CMOSN1323 31 31 D_lateral AREA=3.125E-016    
M1322 45 40 39 45 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1321 39 38 151 45 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1320 38 56 45 45 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1319 45 56 42 45 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1318 42 40 44 45 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1317 42 38 44 45 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1316 31 40 151 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1315 151 38 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1314 38 56 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1313 41 56 44 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1312 44 40 41 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1311 31 38 41 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1310 42 43 45 45 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1309 45 43 40 45 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1308 43 48 45 45 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1307 41 43 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1306 31 43 40 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1305 43 48 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1301 45 46 48 45 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1300 48 117 45 45 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1299 49 117 48 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1298 31 46 49 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1297 are shorted:
* D1297 31 31 D_lateral AREA=3.125E-016    $ (424.5 198 429.5 198.001)CMOSN1297 31 31 D_lateral AREA=3.125E-016    
M1296 59 54 53 59 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1295 53 50 168 59 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1294 50 71 59 59 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1293 59 71 52 59 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1292 52 54 57 59 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1291 52 55 59 59 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1290 52 50 57 59 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1289 31 54 168 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1288 168 50 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1287 50 71 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1286 51 71 57 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1285 51 54 57 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1284 51 55 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1283 31 50 51 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1282 59 55 54 59 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1281 55 62 59 59 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1280 31 55 54 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1279 55 62 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1278 58 117 62 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1277 31 60 58 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1276 are shorted:
* D1276 31 31 D_lateral AREA=3.125E-016    $ (140.5 198 145.5 198.001)CMOSN1276 31 31 D_lateral AREA=3.125E-016    
M1275 59 60 62 59 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1274 62 117 59 59 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1273 74 67 63 74 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1272 63 66 178 74 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1271 31 67 178 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1270 178 66 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1269 66 92 74 74 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1268 74 92 65 74 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1267 65 70 74 74 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1266 74 70 67 74 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1265 65 67 72 74 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1264 65 66 72 74 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1263 66 92 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1262 64 92 72 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1261 64 70 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1260 31 70 67 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1259 64 67 72 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1258 31 66 64 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1257 70 76 74 74 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1256 70 76 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1255 73 117 76 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1254 31 69 73 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1253 are shorted:
* D1253 31 31 D_lateral AREA=3.125E-016    $ (-144 198 -139 198.001)CMOSN1253 31 31 D_lateral AREA=3.125E-016    
M1252 74 69 76 74 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1251 76 117 74 74 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1250 75 191 202 75 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1249 77 84 88 88 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1248 191 200 77 88 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1246 191 84 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1245 31 200 191 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1244 87 203 200 89 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1243 89 206 87 89 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1242 203 103 89 89 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1241 89 103 78 89 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1240 78 206 210 89 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1238 78 203 210 89 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1237 88 90 86 88 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1236 86 79 84 88 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1235 79 85 88 88 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1234 88 85 81 88 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1233 81 90 213 88 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1231 81 79 213 88 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1223 31 90 84 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1222 84 79 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1221 79 85 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1220 80 85 213 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1219 80 90 213 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1217 31 79 80 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1216 88 214 91 88 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1215 89 213 78 89 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M1214 89 213 206 89 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1213 88 91 81 88 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M1212 88 91 90 88 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1211 31 214 91 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1210 93 117 214 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1209 31 95 93 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1206 31 91 80 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M1205 31 91 90 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D1204 are shorted:
* D1204 31 31 D_lateral AREA=3.125E-016    $ (-441 276 -436 276.001)CMOSN1204 31 31 D_lateral AREA=3.125E-016    
M1203 106 100 96 106 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1202 96 99 227 106 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1201 94 95 214 94 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1200 214 117 94 94 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1199 31 100 227 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1198 227 99 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1197 99 119 106 106 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1196 106 119 98 106 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1195 98 104 106 106 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1194 106 104 100 106 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1193 98 100 226 106 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1192 98 99 226 106 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1191 99 119 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1190 97 119 226 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1189 97 104 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1188 31 104 100 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1187 97 100 226 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1186 31 99 97 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1185 104 107 106 106 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1184 106 102 107 106 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1183 104 107 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1182 105 117 107 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1181 31 102 105 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1180 are shorted:
* D1180 31 31 D_lateral AREA=3.125E-016    $ (-725.5 197 -720.5 197.001)CMOSN1180 31 31 D_lateral AREA=3.125E-016    
M1179 106 114 108 106 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1178 108 109 239 106 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1177 107 117 106 106 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1176 31 114 239 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1175 239 109 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1174 109 115 106 106 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1173 106 115 111 106 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1172 111 118 106 106 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1171 106 118 114 106 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1170 111 114 120 106 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1169 111 109 120 106 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1168 109 115 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1167 110 115 120 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1166 110 118 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1165 31 118 114 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1164 110 114 120 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1163 31 109 110 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1162 106 526 118 106 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1161 118 117 106 106 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1160 121 117 118 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1159 31 526 121 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1158 are shorted:
* D1158 31 31 D_lateral AREA=3.125E-016    $ (-1002.5 197 -997.5 197.001)CMOSN1158 31 31 D_lateral AREA=3.125E-016    
* Pins of element D1157 are shorted:
* D1157 31 31 D_lateral AREA=3.125E-016    $ (-1002.5 275 -997.5 275.001)CMOSN1157 31 31 D_lateral AREA=3.125E-016    
M1156 136 245 254 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1155 125 122 135 135 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1154 245 247 125 135 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1153 124 128 247 136 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1152 136 133 124 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1151 135 134 123 135 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1150 123 132 122 135 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1149 31 245 254 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1148 245 122 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1147 31 247 245 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1146 247 128 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1145 31 133 247 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1144 31 134 122 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1143 122 132 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1142 128 44 136 136 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1141 136 44 127 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1140 127 260 136 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1139 136 260 133 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1138 127 133 261 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1137 127 128 261 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1136 132 129 135 135 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1135 135 129 131 135 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1134 131 137 135 135 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1133 135 137 134 135 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1132 131 134 260 135 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1131 131 132 260 135 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1130 128 44 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1129 126 260 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1128 31 260 133 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1127 261 133 126 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1126 31 128 126 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1125 126 44 261 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1124 132 129 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1123 130 129 260 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1122 130 137 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1121 31 137 134 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1120 130 134 260 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1119 31 132 130 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1118 135 262 137 135 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1117 136 33 262 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1116 262 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1115 31 262 137 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1114 138 241 262 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1113 31 33 138 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1112 are shorted:
* D1112 31 31 D_lateral AREA=3.125E-016    $ (696.5 77 701.5 77.001)CMOSN1112 31 31 D_lateral AREA=3.125E-016    
M1111 136 266 282 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1110 142 139 156 156 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1109 266 268 142 156 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1108 141 145 268 136 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1107 136 149 141 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1105 156 150 140 156 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1104 140 148 139 156 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1102 31 266 282 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1101 266 139 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1100 31 268 266 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1099 268 145 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1098 31 149 268 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1096 31 150 139 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1095 139 148 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1093 136 57 145 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M1092 136 57 144 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1091 144 280 136 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1090 136 280 149 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1089 144 149 281 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1088 144 145 281 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1087 156 151 148 156 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M1086 156 151 147 156 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1085 147 153 156 156 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1084 156 153 150 156 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1083 147 150 280 156 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1082 147 148 280 156 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1081 31 57 145 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M1080 143 280 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1079 31 280 149 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1078 281 149 143 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1077 31 145 143 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1076 143 57 281 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1075 31 151 148 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M1074 146 151 280 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1073 146 153 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1072 31 153 150 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1071 146 150 280 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1070 31 148 146 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1069 156 152 153 156 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1068 136 46 152 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1067 152 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1065 157 290 155 173 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1064 31 152 153 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1063 154 241 152 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1062 31 46 154 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1060 31 290 157 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D1059 are shorted:
* D1059 31 31 D_lateral AREA=3.125E-016    $ (412 77 417 77.001)CMOSN1059 31 31 D_lateral AREA=3.125E-016    
M1058 136 157 302 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1057 173 158 155 173 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=562.5f PS=2.25u    
M1056 160 171 290 136 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1055 136 165 160 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1054 171 72 136 136 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1053 136 72 162 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1052 173 166 159 173 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1051 159 170 158 173 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1050 170 168 173 173 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1049 173 168 164 173 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1048 31 157 302 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1047 31 158 157 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=968.75f PS=3u    
M1046 290 171 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1045 31 165 290 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1044 171 72 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1043 31 171 161 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1042 31 166 158 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1041 158 170 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1040 170 168 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1039 31 170 163 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1038 173 172 167 173 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1037 162 299 136 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1036 136 299 165 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1035 162 165 300 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1034 162 171 300 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1033 164 167 173 173 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1032 173 167 166 173 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1031 164 166 299 173 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1030 164 170 299 173 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1029 31 172 167 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1028 169 241 172 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1027 31 60 169 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1026 161 299 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1025 31 299 165 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1024 300 165 161 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M1023 161 72 300 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1022 163 167 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1021 31 167 166 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1020 163 166 299 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1019 163 168 299 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D1018 are shorted:
* D1018 31 31 D_lateral AREA=3.125E-016    $ (128 77 133 77.001)CMOSN1018 31 31 D_lateral AREA=3.125E-016    
M1017 136 60 172 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1016 172 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1015 136 306 313 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1014 174 177 181 181 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1013 306 312 174 181 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1012 31 306 313 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1011 306 177 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1010 31 312 306 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1009 180 175 312 136 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1008 136 186 180 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1007 175 210 136 136 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1006 136 210 183 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1005 183 175 323 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1004 181 187 179 181 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1003 179 176 177 181 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1002 176 178 181 181 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1001 181 178 185 181 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1000 185 176 322 181 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M999 312 175 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M998 31 186 312 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M997 175 210 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M996 31 175 182 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M995 182 210 323 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M994 31 187 177 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M993 177 176 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M992 176 178 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M991 184 178 322 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M990 31 176 184 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M989 181 190 188 181 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M988 183 322 136 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M987 136 322 186 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M986 183 186 323 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M985 185 188 181 181 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M984 181 188 187 181 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M983 185 187 322 181 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M982 31 190 188 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M981 189 241 190 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M980 31 69 189 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M979 182 322 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M978 31 322 186 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M977 323 186 182 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M976 184 188 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M975 31 188 187 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M974 184 187 322 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
* Pins of element D973 are shorted:
* D973 31 31 D_lateral AREA=3.125E-016    $ (-156.5 77 -151.5 77.001)CMOSN973 31 31 D_lateral AREA=3.125E-016    
M972 136 69 190 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M971 190 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M970 136 326 337 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M969 192 201 207 207 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M968 326 336 192 207 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M967 31 191 202 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M966 31 326 337 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M965 326 201 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M964 31 336 326 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M963 205 194 336 136 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M962 136 208 205 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M961 194 226 136 136 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M960 136 226 196 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M959 196 208 343 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M957 196 194 343 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M956 207 209 204 207 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M955 204 197 201 207 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M954 197 202 207 207 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M953 207 202 199 207 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M952 199 209 342 207 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M950 199 197 342 207 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M949 200 206 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M948 200 203 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M947 31 103 203 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M946 193 103 210 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M945 31 203 193 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M944 193 206 210 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M942 336 194 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M941 31 208 336 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M940 194 226 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M939 343 208 195 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M937 31 194 195 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M936 195 226 343 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M935 31 209 201 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M934 201 197 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M933 197 202 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M932 198 202 342 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M931 198 209 342 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M929 31 197 198 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M928 207 215 211 207 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M927 136 342 196 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M926 136 342 208 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M925 207 211 199 207 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M924 207 211 209 207 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M923 31 213 206 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M922 31 213 193 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M921 31 215 211 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M920 212 241 215 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M919 31 95 212 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M918 31 342 195 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M917 31 342 208 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M916 31 211 198 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M915 31 211 209 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D914 are shorted:
* D914 31 31 D_lateral AREA=3.125E-016    $ (-441 173 -436 173.001)CMOSN914 31 31 D_lateral AREA=3.125E-016    
* Pins of element D913 are shorted:
* D913 31 31 D_lateral AREA=3.125E-016    $ (-441 77 -436 77.001)CMOSN913 31 31 D_lateral AREA=3.125E-016    
M912 136 95 215 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M911 215 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M910 136 346 359 136 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M909 218 225 228 228 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M908 346 358 218 228 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M906 136 229 217 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M905 228 230 216 228 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M903 31 346 359 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M902 346 225 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M901 31 358 346 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M900 31 229 358 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M899 31 230 225 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M898 358 219 217 136 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M897 219 120 136 136 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M896 136 120 221 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M895 221 229 363 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M894 221 362 136 136 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M893 136 362 229 136 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M892 221 219 363 136 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M891 225 222 216 228 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M890 222 227 228 228 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M889 228 227 224 228 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M888 224 230 362 228 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M887 224 231 228 228 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M886 228 231 230 228 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M885 224 222 362 228 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M884 358 219 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M883 219 120 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M882 363 229 220 31 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M881 220 362 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M880 31 362 229 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M879 31 219 220 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M878 220 120 363 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M877 225 222 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M876 222 227 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M875 223 227 362 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M874 223 230 362 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M873 223 231 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M872 31 231 230 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M871 31 222 223 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M870 228 233 231 228 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M869 136 102 233 136 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M868 31 233 231 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M867 232 241 233 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M866 31 102 232 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D865 are shorted:
* D865 31 31 D_lateral AREA=3.125E-016    $ (-725.5 77 -720.5 77.001)CMOSN865 31 31 D_lateral AREA=3.125E-016    
M864 240 238 234 240 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M863 234 235 372 240 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M862 233 241 136 136 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M861 31 238 372 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M860 372 235 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M859 235 239 240 240 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M858 240 239 237 240 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M857 237 242 240 240 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M856 240 242 238 240 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M855 237 238 243 240 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M854 237 235 243 240 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M853 235 239 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M852 236 239 243 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M851 236 242 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M850 31 242 238 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M849 236 238 243 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M848 31 235 236 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M847 240 526 242 240 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M846 242 241 240 240 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M845 244 241 242 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M844 31 526 244 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D843 are shorted:
* D843 31 31 D_lateral AREA=3.125E-016    $ (-1002.5 102 -997.5 102.001)CMOSN843 31 31 D_lateral AREA=3.125E-016    
M842 263 381 396 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M841 250 246 287 287 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M840 381 382 250 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M839 263 258 249 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M838 249 253 382 263 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M837 287 259 248 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M836 248 257 246 287 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M835 31 381 396 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M834 381 246 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M833 31 382 381 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M832 31 258 382 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M831 382 253 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M830 31 259 246 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M829 246 257 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M828 253 281 263 263 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M827 263 281 252 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M826 252 394 263 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M825 263 394 258 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M824 252 258 395 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M823 252 253 395 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M822 257 254 287 287 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M821 287 254 256 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M820 256 264 287 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M819 287 264 259 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M818 256 259 394 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M817 256 257 394 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M816 253 281 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M815 251 281 395 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M814 251 394 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M813 31 394 258 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M812 251 258 395 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M811 31 253 251 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M810 257 254 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M809 255 254 394 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M808 255 264 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M807 31 264 259 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M806 255 259 394 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M805 31 257 255 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M804 287 398 264 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M803 263 33 398 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M802 398 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M801 31 398 264 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M800 265 374 398 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M799 31 33 265 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D798 are shorted:
* D798 31 31 D_lateral AREA=3.125E-016    $ (696.5 -19 701.5 -18.999)CMOSN798 31 31 D_lateral AREA=3.125E-016    
M797 263 407 424 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M796 271 267 287 287 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M795 407 408 271 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M794 263 278 270 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M793 270 274 408 263 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M791 287 279 269 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M790 269 277 267 287 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M788 31 407 424 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M787 407 267 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M786 31 408 407 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M785 31 278 408 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M784 408 274 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M782 31 279 267 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M781 267 277 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M779 263 300 274 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M778 263 300 273 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M777 273 421 263 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M776 263 421 278 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M775 273 278 422 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M774 273 274 422 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M773 287 282 277 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M772 287 282 276 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M771 276 284 287 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M770 287 284 279 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M769 276 279 421 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M768 276 277 421 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M767 31 300 274 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M766 272 300 422 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M765 272 421 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M764 31 421 278 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M763 272 278 422 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M762 31 274 272 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M761 31 282 277 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M760 275 282 421 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M759 275 284 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M758 31 284 279 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M757 275 279 421 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M756 31 277 275 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M755 287 283 284 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M754 263 46 283 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M753 283 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M751 288 430 286 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M750 31 283 284 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M749 285 374 283 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M748 31 46 285 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M746 31 430 288 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D745 are shorted:
* D745 31 31 D_lateral AREA=3.125E-016    $ (412 -19 417 -18.999)CMOSN745 31 31 D_lateral AREA=3.125E-016    
M744 263 288 446 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M743 287 289 286 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=562.5f PS=2.25u    
M742 263 297 292 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M741 292 305 430 263 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M740 305 323 263 263 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M739 263 323 294 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M738 287 298 291 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M737 291 304 289 287 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M736 304 302 287 287 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M735 287 302 296 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M734 31 288 446 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M733 31 289 288 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=968.75f PS=3u    
M732 31 297 430 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M731 430 305 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M730 305 323 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M729 31 305 293 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M728 31 298 289 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M727 289 304 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M726 304 302 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M725 31 304 295 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M724 287 307 301 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M723 294 443 263 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M722 263 443 297 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M721 294 297 444 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M720 294 305 444 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M719 296 301 287 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M718 287 301 298 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M717 296 298 443 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M716 296 304 443 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M715 31 307 301 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M714 303 374 307 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M713 31 60 303 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M712 293 443 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M711 31 443 297 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M710 293 297 444 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M709 293 323 444 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M708 295 301 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M707 31 301 298 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M706 295 298 443 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M705 295 302 443 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D704 are shorted:
* D704 31 31 D_lateral AREA=3.125E-016    $ (128 -19 133 -18.999)CMOSN704 31 31 D_lateral AREA=3.125E-016    
M703 263 60 307 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M702 307 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M701 263 450 464 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M700 308 311 287 287 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M699 450 454 308 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M698 31 450 464 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M697 450 311 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M696 31 454 450 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M695 263 320 315 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M694 315 309 454 263 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M693 309 343 263 263 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M692 263 343 317 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M691 317 309 461 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M690 287 321 314 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M689 314 310 311 287 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M688 310 313 287 287 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M687 287 313 319 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M686 319 310 460 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M685 31 320 454 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M684 454 309 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M683 309 343 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M682 316 343 461 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M681 31 309 316 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M680 31 321 311 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M679 311 310 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M678 310 313 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M677 318 313 460 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M676 31 310 318 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M675 287 327 324 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M674 317 460 263 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M673 263 460 320 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M672 317 320 461 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M671 319 324 287 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M670 287 324 321 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M669 319 321 460 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M668 31 327 324 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M667 325 374 327 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M666 31 69 325 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M665 316 460 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M664 31 460 320 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M663 316 320 461 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M662 318 324 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M661 31 324 321 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M660 318 321 460 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
* Pins of element D659 are shorted:
* D659 31 31 D_lateral AREA=3.125E-016    $ (-156.5 -19 -151.5 -18.999)CMOSN659 31 31 D_lateral AREA=3.125E-016    
M658 263 69 327 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M657 327 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M656 263 473 480 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M655 328 335 287 287 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M654 473 479 328 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M653 31 473 480 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M652 473 335 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M651 31 479 473 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M650 263 340 339 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M649 339 329 479 263 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M648 329 363 263 263 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M647 263 363 331 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M646 331 340 489 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M644 331 329 489 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M643 287 341 338 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M642 338 332 335 287 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M641 332 337 287 287 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M640 287 337 334 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M639 334 341 488 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M637 334 332 488 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M636 31 340 479 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M635 479 329 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M634 329 363 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M633 330 363 489 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M632 330 340 489 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M630 31 329 330 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M629 31 341 335 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M628 335 332 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M627 332 337 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M626 333 337 488 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M625 333 341 488 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M623 31 332 333 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M622 287 347 344 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M621 263 488 331 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M620 263 488 340 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M619 287 344 334 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M618 287 344 341 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M617 31 347 344 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M616 345 374 347 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M615 31 95 345 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M614 31 488 330 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M613 31 488 340 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M612 31 344 333 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M611 31 344 341 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D610 are shorted:
* D610 31 31 D_lateral AREA=3.125E-016    $ (-441 -19 -436 -18.999)CMOSN610 31 31 D_lateral AREA=3.125E-016    
M609 263 95 347 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M608 347 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M607 263 496 507 263 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M606 350 357 287 287 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M605 496 506 350 287 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M604 263 360 349 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M602 287 361 348 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M600 31 496 507 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M599 496 357 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M598 31 506 496 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M597 31 360 506 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M596 31 361 357 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M595 506 351 349 263 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M594 351 243 263 263 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M593 263 243 353 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M592 353 360 514 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M591 353 513 263 263 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M590 263 513 360 263 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M589 353 351 514 263 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M588 357 354 348 287 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M587 354 359 287 287 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M586 287 359 356 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M585 356 361 513 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M584 356 364 287 287 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M583 287 364 361 287 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M582 356 354 513 287 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M581 506 351 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M580 351 243 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M579 352 243 514 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M578 352 360 514 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M577 352 513 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M576 31 513 360 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M575 31 351 352 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M574 357 354 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M573 354 359 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M572 355 359 513 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M571 355 361 513 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M570 355 364 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M569 31 364 361 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M568 31 354 355 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M567 287 366 364 287 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M566 263 102 366 263 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M565 31 366 364 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M564 365 374 366 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M563 31 102 365 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D562 are shorted:
* D562 31 31 D_lateral AREA=3.125E-016    $ (-725.5 -19 -720.5 -18.999)CMOSN562 31 31 D_lateral AREA=3.125E-016    
M561 373 371 367 373 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M560 367 368 524 373 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M559 366 374 263 263 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M558 31 371 524 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M557 524 368 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M556 368 372 373 373 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M555 373 372 370 373 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M554 370 375 373 373 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M553 373 375 371 373 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M552 370 371 376 373 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M551 370 368 376 373 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M550 368 372 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M549 369 372 376 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M548 369 375 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M547 31 375 371 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M546 369 371 376 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M545 31 368 369 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M544 373 526 375 373 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M543 375 374 373 373 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M542 377 374 375 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M541 31 526 377 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D540 are shorted:
* D540 31 31 D_lateral AREA=3.125E-016    $ (-1002.5 6 -997.5 6.001)CMOSN540 31 31 D_lateral AREA=3.125E-016    
M539 399 378 536 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M538 385 379 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M537 378 380 385 400 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M536 399 392 384 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M535 384 386 380 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M534 400 393 383 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M533 383 389 379 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M532 31 378 536 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M531 378 379 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M530 31 380 378 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M529 31 392 380 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M528 380 386 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M527 31 393 379 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M526 379 389 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M525 386 422 399 399 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M524 399 422 388 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M523 388 397 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M522 399 397 392 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M521 388 392 402 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M520 388 386 402 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M519 389 396 400 400 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M518 400 396 391 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M517 391 401 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M516 400 401 393 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M515 391 393 397 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M514 391 389 397 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M513 386 422 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M512 387 422 402 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M511 387 397 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M510 31 397 392 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M509 387 392 402 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M508 31 386 387 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M507 389 396 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M506 390 396 397 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M505 390 401 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M504 31 401 393 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M503 390 393 397 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M502 31 389 390 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M501 400 33 401 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M500 401 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M499 403 528 401 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M498 31 33 403 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D497 are shorted:
* D497 31 31 D_lateral AREA=3.125E-016    $ (696.5 -64 701.5 -63.999)CMOSN497 31 31 D_lateral AREA=3.125E-016    
M496 399 404 556 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M495 411 405 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M494 404 406 411 400 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M493 399 418 410 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M492 410 414 406 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M491 400 420 409 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M490 409 417 405 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M489 31 404 556 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M488 404 405 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M487 31 406 404 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M486 31 418 406 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M485 406 414 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M484 31 420 405 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M483 405 417 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M482 414 444 399 399 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M481 399 444 413 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M480 413 419 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M479 399 419 418 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M478 413 418 423 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M477 413 414 423 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M476 417 424 400 400 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M475 400 424 416 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M474 416 425 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M473 400 425 420 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M472 416 420 419 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M471 416 417 419 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M470 414 444 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M469 412 444 423 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M468 412 419 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M467 31 419 418 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M466 412 418 423 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M465 31 414 412 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M464 417 424 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M463 415 424 419 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M462 415 425 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M461 31 425 420 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M460 415 420 419 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M459 31 417 415 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M457 400 46 425 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M456 425 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M454 426 528 425 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M453 31 46 426 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D452 are shorted:
* D452 31 31 D_lateral AREA=3.125E-016    $ (412 -64 417 -63.999)CMOSN452 31 31 D_lateral AREA=3.125E-016    
M451 399 427 574 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M450 433 428 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M449 433 429 427 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=2.3125p PS=7u    
M448 399 440 432 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M447 432 436 429 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M446 399 461 436 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M445 400 442 431 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M444 431 439 428 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M443 400 446 439 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M442 31 427 574 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M441 427 428 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M440 427 429 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.9375p PS=6u    
M439 31 440 429 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M438 429 436 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M437 31 461 436 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M436 31 442 428 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M435 428 439 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M434 31 446 439 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M433 435 441 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M432 399 441 440 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M431 435 440 445 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M430 435 436 445 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M429 399 461 435 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M428 438 449 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M427 400 449 442 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M426 438 442 441 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M425 438 439 441 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M424 400 446 438 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M423 447 528 449 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M422 31 60 447 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M421 434 441 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M420 31 441 440 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M419 434 440 445 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M418 31 436 434 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M417 434 461 445 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M416 437 449 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M415 31 449 442 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M414 437 442 441 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M413 31 439 437 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M412 437 446 441 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D411 are shorted:
* D411 31 31 D_lateral AREA=3.125E-016    $ (128 -64 133 -63.999)CMOSN411 31 31 D_lateral AREA=3.125E-016    
M410 399 448 587 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M409 451 452 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M408 448 453 451 400 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M407 400 60 449 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M406 449 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M405 31 448 587 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M404 448 452 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M403 31 453 448 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M402 399 457 456 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M401 456 470 453 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M400 470 489 399 399 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M399 399 489 469 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M398 400 459 455 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M397 455 468 452 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M396 468 464 400 400 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M395 400 464 467 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M394 31 457 453 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M393 453 470 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M392 470 489 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M391 31 470 465 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M390 31 459 452 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M389 452 468 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M388 468 464 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M387 31 468 463 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M386 469 458 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M385 399 458 457 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M384 469 457 462 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M383 469 470 462 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M382 467 472 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M381 400 472 459 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M380 467 459 458 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M379 467 468 458 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M378 466 528 472 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M377 31 69 466 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M376 465 458 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M375 31 458 457 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M374 465 457 462 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M373 465 489 462 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M372 463 472 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M371 31 472 459 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M370 463 459 458 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M369 463 464 458 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D368 are shorted:
* D368 31 31 D_lateral AREA=3.125E-016    $ (-156.5 -64 -151.5 -63.999)CMOSN368 31 31 D_lateral AREA=3.125E-016    
M367 399 471 600 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M366 474 478 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M365 471 477 474 400 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M364 400 69 472 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M363 472 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M362 31 471 600 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M361 471 478 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M360 31 477 471 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M359 399 493 482 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M358 482 475 477 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M357 475 514 399 399 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M356 399 514 484 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M354 484 475 490 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M353 400 492 481 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M352 481 476 478 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M351 476 480 400 400 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M350 400 480 486 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M348 486 476 487 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M347 31 493 477 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M346 477 475 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M345 475 514 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M344 483 514 490 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M342 31 475 483 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M341 31 492 478 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M340 478 476 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M339 476 480 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M338 485 480 487 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M336 31 476 485 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M335 484 487 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M334 399 487 493 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M333 484 493 490 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M332 486 495 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M331 400 495 492 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M330 486 492 487 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M329 491 528 495 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M328 31 95 491 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M327 483 487 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M326 31 487 493 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M325 483 493 490 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M324 485 495 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M323 31 495 492 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M322 485 492 487 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
* Pins of element D321 are shorted:
* D321 31 31 D_lateral AREA=3.125E-016    $ (-441 -64 -436 -63.999)CMOSN321 31 31 D_lateral AREA=3.125E-016    
M320 399 494 622 399 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M319 497 505 400 400 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M318 494 504 497 400 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M317 400 95 495 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M316 495 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M315 31 494 622 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M314 494 505 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M313 31 504 494 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M312 399 510 509 399 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M311 509 498 504 399 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M310 498 376 399 399 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M309 399 376 500 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M308 500 510 515 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M307 500 512 399 399 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M306 500 498 515 399 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M305 400 511 508 400 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M304 508 501 505 400 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M303 501 507 400 400 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M302 400 507 503 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M301 503 511 512 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M300 503 518 400 400 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M299 503 501 512 400 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M298 31 510 504 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M297 504 498 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M296 498 376 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M295 499 376 515 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M294 499 510 515 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M293 499 512 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M292 31 498 499 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M291 31 511 505 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M290 505 501 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M289 501 507 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M288 502 507 512 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M287 502 511 512 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M286 502 518 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M285 31 501 502 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M284 400 102 518 400 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M283 399 512 510 399 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M282 400 518 511 400 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M281 516 528 518 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M280 31 102 516 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M279 31 512 510 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M278 31 518 511 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D277 are shorted:
* D277 31 31 D_lateral AREA=3.125E-016    $ (-725.5 -64 -720.5 -63.999)CMOSN277 31 31 D_lateral AREA=3.125E-016    
M276 518 528 400 400 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M275 527 521 517 527 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M274 517 525 640 527 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M273 527 524 525 527 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M271 31 521 640 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M270 640 525 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M269 31 524 525 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M267 520 522 527 527 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M266 527 522 521 527 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M265 520 521 523 527 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M264 520 525 523 527 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M263 520 524 527 527 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M262 522 529 527 527 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M261 519 522 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M260 31 522 521 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M259 519 521 523 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M258 519 525 31 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M257 519 524 523 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M256 522 529 31 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M255 527 526 529 527 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M254 529 528 527 527 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M253 530 528 529 31 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M252 31 526 530 31 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D251 are shorted:
* D251 31 31 D_lateral AREA=3.125E-016    $ (-1002.5 -89 -997.5 -88.999)CMOSN251 31 31 D_lateral AREA=3.125E-016    
M250 537 535 531 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M249 531 532 555 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M248 31 535 555 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M247 555 532 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M246 532 536 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M245 537 536 534 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M244 534 423 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M243 537 423 535 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M242 534 535 538 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M241 534 532 538 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M240 532 536 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M239 533 536 538 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M238 533 423 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M237 31 423 535 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M236 533 535 538 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M235 31 532 533 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M234 557 539 575 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M233 544 540 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M232 539 541 544 537 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M231 557 551 543 557 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M230 543 547 541 557 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M229 537 554 542 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M228 542 550 540 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M227 31 539 575 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M226 539 540 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M225 31 541 539 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M224 31 551 541 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M223 541 547 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M222 31 554 540 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M221 540 550 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M220 547 555 557 557 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M219 557 555 546 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M218 546 552 557 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M217 557 552 551 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M216 546 551 553 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M215 546 547 553 557 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M214 550 556 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M213 537 556 549 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M212 549 445 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M211 537 445 554 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M210 549 554 552 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M209 549 550 552 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M208 547 555 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M207 545 555 553 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M206 545 552 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M205 31 552 551 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M204 545 551 553 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M203 31 547 545 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M202 550 556 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M201 548 556 552 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M200 548 445 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M199 31 445 554 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M198 548 554 552 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M197 31 550 548 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M194 557 558 589 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M193 563 559 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M192 563 560 558 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=2.3125p PS=7u    
M191 557 570 562 557 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M190 562 566 560 557 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M189 557 575 566 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M188 537 573 561 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M187 561 569 559 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M186 537 574 569 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M185 31 558 589 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M184 558 559 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M183 558 560 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.9375p PS=6u    
M182 31 570 560 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M181 560 566 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M180 31 575 566 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M179 31 573 559 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M178 559 569 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M177 31 574 569 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M176 565 571 557 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M175 557 571 570 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M174 565 570 572 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M173 565 566 572 557 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M172 557 575 565 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M171 568 462 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M170 537 462 573 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M169 568 573 571 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M168 568 569 571 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M167 537 574 568 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M166 564 571 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M165 31 571 570 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M164 564 570 572 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M163 31 566 564 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M162 564 575 572 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M161 567 462 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M160 31 462 573 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M159 567 573 571 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M158 31 569 567 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M157 567 574 571 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M156 557 576 609 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M155 577 578 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M154 576 579 577 537 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M153 31 576 609 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M152 576 578 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M151 31 579 576 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M150 557 582 581 557 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M149 581 593 579 557 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M148 593 589 557 557 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M147 557 589 592 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M146 537 585 580 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M145 580 591 578 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M144 591 587 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M143 537 587 590 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M142 31 582 579 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M141 579 593 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M140 593 589 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M139 31 593 588 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M138 31 585 578 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M137 578 591 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M136 591 587 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M135 31 591 586 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M134 592 583 557 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M133 557 583 582 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M132 592 582 584 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M131 592 593 584 557 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M130 590 490 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M129 537 490 585 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M128 590 585 583 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M127 590 591 583 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M126 588 583 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M125 31 583 582 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M124 588 582 584 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M123 588 589 584 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M122 586 490 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M121 31 490 585 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M120 586 585 583 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M119 586 587 583 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M118 557 594 629 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M117 595 599 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M116 594 598 595 537 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M115 31 594 629 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M114 594 599 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M113 31 598 594 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M112 557 611 602 557 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M111 602 596 598 557 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M110 596 609 557 557 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M109 557 609 604 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M107 604 596 608 557 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M106 537 610 601 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M105 601 597 599 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M104 597 600 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M103 537 600 606 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M101 606 597 607 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M100 31 611 598 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M99 598 596 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M98 596 609 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M97 603 609 608 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M95 31 596 603 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M94 31 610 599 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M93 599 597 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M92 597 600 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M91 605 600 607 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M89 31 597 605 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M88 604 607 557 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M87 557 607 611 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M86 604 611 608 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M85 606 515 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M84 537 515 610 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M83 606 610 607 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M82 603 607 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M81 31 607 611 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M80 603 611 608 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M79 605 515 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M78 31 515 610 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M77 605 610 607 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M76 557 612 642 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M75 613 621 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M74 612 620 613 537 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M73 31 612 642 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M72 612 621 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M71 31 620 612 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M70 557 625 624 557 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M69 624 614 620 557 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M68 614 629 557 557 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M67 557 629 616 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M66 616 625 628 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M65 616 627 557 557 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M64 616 614 628 557 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M63 537 626 623 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M62 623 617 621 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M61 617 622 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M60 537 622 619 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M59 619 626 627 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M58 619 523 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M57 619 617 627 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M56 31 625 620 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M55 620 614 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M54 614 629 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M53 615 629 628 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M52 615 625 628 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M51 615 627 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M50 31 614 615 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M49 31 626 621 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M48 621 617 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M47 617 622 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M46 618 622 627 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M45 618 626 627 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M44 618 523 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M43 31 617 618 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M42 557 627 625 557 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M41 537 523 626 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M40 31 627 625 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M39 31 523 626 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M38 557 630 631 557 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M37 632 641 537 537 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M36 630 639 632 537 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M35 31 630 631 31 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M34 630 641 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M33 31 639 630 31 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M32 649 645 644 649 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M31 644 633 639 649 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M30 633 640 649 649 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M29 649 640 635 649 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M28 635 645 648 649 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M27 635 647 649 649 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M26 635 633 648 649 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M25 537 646 643 537 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M24 643 636 641 537 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M23 636 642 537 537 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M22 537 642 638 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M21 638 646 647 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M20 638 537 537 537 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M19 638 636 647 537 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M18 31 645 639 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M17 639 633 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M16 633 640 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M15 634 640 648 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M14 634 645 648 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M13 634 647 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M12 31 633 634 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M11 31 646 641 31 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M10 641 636 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M9 636 642 31 31 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M8 637 642 647 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M7 637 646 647 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M6 637 537 31 31 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M5 31 636 637 31 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M4 649 647 645 649 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3 537 537 646 537 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2 31 647 645 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1 31 537 646 31 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    

* Total Nodes: 649
* Total Elements: 1367
* Total Number of Shorted Elements not written to the SPICE file: 0
* Output Generation Elapsed Time: 0.047 sec
* Total Extract Elapsed Time: 1.797 sec

* INPUTS 

v1 1 0 5v
v2 3 0 5v
v3 7 0 5v
v4 10 0 5v
v5 16 0 5v
v6 22 0 5v
v7 32 0 5v
v8 45 0 5v
v9 59 0 5v
v10 74 0 5v
v11 75 0 5v 
v12 88 0 5v
v13 89 0 5v
v14 94 0 5v
v15 106 0 5v
v16 135 0 5v
v17 136 0 5v
v18 156 0 5v 
v19 173 0 5v
v20 181 0 5v
v21 207 0 5v
v22 228 0 5v
v23 240 0 5v
v24 263 0 5v
v25 287 0 5v
v26 373 0 5v
v27 399 0 5v
v28 400 0 5v
v29 527 0 5v
v30 537 0 5v
v31 557 0 5v
v32 649 0 5v
v33 31 0 0v


v34 9 0 pulse(0 5v 50n 0.05n 0.05n 250n 100n)
v35 117 0 0v
v36 241 0 0v
v37 374 0 0v
v38 528 0 0v

v39 33 0 5v
v40 46 0 5v
v41 60 0 5v
v42 69 0 5v
v43 95 0 5v
v44 102 0 5v
v45 526 0 pulse(0v 5v 50n 0.05n 0.05n 250n 100n)
* OUTPUTS 
* OUTPUT can be put in trace in simulation 
* 
.op
.tran 0.1ns 200ns
.probe
.END