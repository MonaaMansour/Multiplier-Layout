
* Circuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 ;CMOSNuit Extracted by Tanner Research's L-Edit Version 15.00 / Extract Version 15.00 
* TDB File:  C:\Documents and Settings\Owner\Desktop\Project\Multiplier_pads.tdb
* Cell:  Cell0	Version 1.12
* Extract Definition File:  ..\extract\mhp_n05.ext
* Extract Date and Time:  01/31/2023 - 01:32

* Tech: AMI_C5N
* LOT: T22Y_TT (typical)                  WAF: 3104
* Temperature_parameters=Optimized 
.MODEL CMOSN NMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6696061
+K1      = 0.8351612      K2      = -0.0839158     K3      = 23.1023856
+K3B     = -7.6841108     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.9047241      DVT1    = 0.4302695      DVT2    = -0.134857
+U0      = 458.439679     UA      = 1E-13          UB      = 1.485499E-18
+UC      = 1.629939E-11   VSAT    = 1.643993E5     A0      = 0.6103537
+AGS     = 0.1194608      B0      = 2.674756E-6    B1      = 5E-6
+KETA    = -2.640681E-3   A1      = 8.219585E-5    A2      = 0.3564792
+RDSW    = 1.387108E3     PRWG    = 0.0299916      PRWB    = 0.0363981
+WR      = 1              WINT    = 2.472348E-7    LINT    = 3.597605E-8
+XL      = 0              XW      = 0              DWG     = -1.287163E-8
+DWB     = 5.306586E-8    VOFF    = 0              NFACTOR = 0.8365585
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.0246738      ETAB    = -1.406123E-3
+DSUB    = 0.2543458      PCLM    = 2.5945188      PDIBLC1 = -0.4282336
+PDIBLC2 = 2.311743E-3    PDIBLCB = -0.0272914     DROUT   = 0.7283566
+PSCBE1  = 5.598623E8     PSCBE2  = 5.461645E-5    PVAG    = 0
+DELTA   = 0.01           RSH     = 81.8           MOBMOD  = 1
+PRT     = 8.621          UTE     = -1             KT1     = -0.2501
+KT1L    = -2.58E-9       KT2     = 0              UA1     = 5.4E-10
+UB1     = -4.8E-19       UC1     = -7.5E-11       AT      = 1E5
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2E-10          CGSO    = 2E-10          CGBO    = 1E-9
+CJ      = 4.197772E-4    PB      = 0.99           MJ      = 0.4515044
+CJSW    = 3.242724E-10   PBSW    = 0.1            MJSW    = 0.1153991
+CJSWG   = 1.64E-10       PBSWG   = 0.1            MJSWG   = 0.1153991
+CF      = 0              PVTH0   = 0.0585501      PRDSW   = 133.285505
+PK2     = -0.0299638     WKETA   = -0.0248758     LKETA   = 1.173187E-3
+AF      = 1              KF      = 0)
*
.MODEL CMOSP PMOS (                                LEVEL   = 7
+VERSION = 3.1            TNOM    = 27             TOX     = 1.39E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9214347
+K1      = 0.5553722      K2      = 8.763328E-3    K3      = 6.3063558
+K3B     = -0.6487362     W0      = 1.280703E-8    NLX     = 2.593997E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 2.5131165      DVT1    = 0.5480536      DVT2    = -0.1186489
+U0      = 212.0166131    UA      = 2.807115E-9    UB      = 1E-21
+UC      = -5.82128E-11   VSAT    = 1.713601E5     A0      = 0.8430019
+AGS     = 0.1328608      B0      = 7.117912E-7    B1      = 5E-6
+KETA    = -3.674859E-3   A1      = 4.77502E-5     A2      = 0.3
+RDSW    = 2.837206E3     PRWG    = -0.0363908     PRWB    = -1.016722E-5
+WR      = 1              WINT    = 2.838038E-7    LINT    = 5.528807E-8
+XL      = 0              XW      = 0              DWG     = -1.606385E-8
+DWB     = 2.266386E-8    VOFF    = -0.0558512     NFACTOR = 0.9342488
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.3251882      ETAB    = -0.0580325
+DSUB    = 1              PCLM    = 2.2409567      PDIBLC1 = 0.0411445
+PDIBLC2 = 3.355575E-3    PDIBLCB = -0.0551797     DROUT   = 0.2036901
+PSCBE1  = 6.44809E9      PSCBE2  = 6.300848E-10   PVAG    = 0
+DELTA   = 0.01           RSH     = 101.6          MOBMOD  = 1
+PRT     = 59.494         UTE     = -1             KT1     = -0.2942
+KT1L    = 1.68E-9        KT2     = 0              UA1     = 4.5E-9
+UB1     = -6.3E-18       UC1     = -1E-10         AT      = 1E3
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.9E-10        CGSO    = 2.9E-10        CGBO    = 1E-9
+CJ      = 7.235528E-4    PB      = 0.9527355      MJ      = 0.4955293
+CJSW    = 2.692786E-10   PBSW    = 0.99           MJSW    = 0.2958392
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.2958392
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 5.292165E-3    LKETA   = -4.205905E-3 
+AF      = 1              KF      = 0)
*

* Warning:  Layers with Unassigned AREA Capacitance.
*   <n well wire>
*   <subs>
*   <allsubs>
*   <poly wire>
*   <Metal1>
*   <Metal1-Tight>
*   <Metal2>
*   <Metal2-Tight>
*   <LPNP emitter>
*   <LPNP collector>
* Warning:  Layers with Unassigned FRINGE Capacitance.
*   <Pad Comment>
*   <ndiff>
*   <n well wire>
*   <pdiff>
*   <subs>
*   <allsubs>
*   <AllMetal1>
*   <poly wire>
*   <AllMetal2>
*   <Metal3>
*   <Metal1>
*   <Metal1-Tight>
*   <Metal2>
*   <Metal2-Tight>
*   <LPNP emitter>
*   <LPNP collector>

* NODE NAME ALIASES
*       1 = U320/DataInUnBuf (1221.5 , 446)
*       2 = U319/DataInUnBuf (785.5 , 446)
*       3 = U318/DataInUnBuf (349.5 , 446)
*       4 = U317/DataInUnBuf (-86.5 , 446)
*       5 = U316/DataInUnBuf (-522.5 , 446)
*       6 = U315/DataInUnBuf (-958.5 , 446)
*       7 = U313/DataInUnBuf (-1394.5 , 446)
*       8 = U310/U228/VDD (-716 , -933.5)
*       8 = U331/VddWell (-1557.5 , -2302)
*       8 = U330/VddWell (-1557.5 , -2302)
*       8 = U331/VddSel (-1557.5 , -2301)
*       8 = U331/VddAct (-1557.5 , -2299)
*       8 = U330/VddSel (-1557.5 , -2301)
*       8 = U330/VddAct (-1557.5 , -2299)
*       8 = U331/Vdd (-1557.5 , -2234)
*       8 = U331/Vdd2 (-1557.5 , -2299)
*       8 = U330/Vdd (-1557.5 , -2234)
*       8 = U330/Vdd2 (-1557.5 , -2299)
*       8 = U332/VddWell (-1121.5 , -2302)
*       8 = U332/VddSel (-1121.5 , -2301)
*       8 = U332/VddAct (-1121.5 , -2299)
*       8 = U332/Vdd (-1121.5 , -2234)
*       8 = U332/Vdd2 (-1121.5 , -2299)
*       8 = U333/VddWell (-685.5 , -2302)
*       8 = U333/VddSel (-685.5 , -2301)
*       8 = U333/VddAct (-685.5 , -2299)
*       8 = U333/Vdd (-685.5 , -2234)
*       8 = U333/Vdd2 (-685.5 , -2299)
*       8 = U334/VddWell (-249.5 , -2302)
*       8 = U334/VddSel (-249.5 , -2301)
*       8 = U334/VddAct (-249.5 , -2299)
*       8 = U334/Vdd (-249.5 , -2234)
*       8 = U334/Vdd2 (-249.5 , -2299)
*       8 = U335/VddWell (186.5 , -2302)
*       8 = U335/VddSel (186.5 , -2301)
*       8 = U335/VddAct (186.5 , -2299)
*       8 = U335/Vdd (186.5 , -2234)
*       8 = U335/Vdd2 (186.5 , -2299)
*       8 = U336/VddWell (622.5 , -2302)
*       8 = U336/VddSel (622.5 , -2301)
*       8 = U336/VddAct (622.5 , -2299)
*       8 = U336/Vdd (622.5 , -2234)
*       8 = U336/Vdd2 (622.5 , -2299)
*       8 = U337/VddWell (1058.5 , -2302)
*       8 = U337/VddSel (1058.5 , -2301)
*       8 = U337/VddAct (1058.5 , -2299)
*       8 = U337/Vdd (1058.5 , -2234)
*       8 = U337/Vdd2 (1058.5 , -2299)
*       8 = U338/VddWell (1494.5 , -2302)
*       8 = U338/VddSel (1494.5 , -2301)
*       8 = U338/VddAct (1494.5 , -2299)
*       8 = U338/Vdd (1494.5 , -2234)
*       8 = U338/Vdd2 (1494.5 , -2299)
*       8 = U344/VddWell (-1685.5 , -2170)
*       8 = U344/VddSel (-1684.5 , -2170)
*       8 = U344/VddAct (-1682.5 , -2170)
*       8 = U344/Vdd (-1617.5 , -2170)
*       8 = U344/Vdd2 (-1682.5 , -2170)
*       8 = U339/VddWell (1491.5 , -2174)
*       8 = U339/VddSel (1492.5 , -2174)
*       8 = U339/VddAct (1494.5 , -2174)
*       8 = U339/Vdd (1494.5 , -2174)
*       8 = U339/Vdd2 (1559.5 , -2174)
*       8 = U324/VddWell (-1685.5 , -1734)
*       8 = U324/VddSel (-1684.5 , -1734)
*       8 = U324/VddAct (-1682.5 , -1734)
*       8 = U324/Vdd (-1617.5 , -1734)
*       8 = U324/Vdd2 (-1682.5 , -1734)
*       8 = U340/VddWell (1491.5 , -1738)
*       8 = U340/VddSel (1492.5 , -1738)
*       8 = U340/VddAct (1494.5 , -1738)
*       8 = U340/Vdd (1494.5 , -1738)
*       8 = U340/Vdd2 (1559.5 , -1738)
*       8 = U325/VddWell (-1685.5 , -1298)
*       8 = U325/VddSel (-1684.5 , -1298)
*       8 = U325/VddAct (-1682.5 , -1298)
*       8 = U325/Vdd (-1617.5 , -1298)
*       8 = U325/Vdd2 (-1682.5 , -1298)
*       8 = U341/VddWell (1491.5 , -1302)
*       8 = U341/VddSel (1492.5 , -1302)
*       8 = U341/VddAct (1494.5 , -1302)
*       8 = U341/Vdd (1494.5 , -1302)
*       8 = U341/Vdd2 (1559.5 , -1302)
*       8 = U303/U210/B (-989 , -1041.5)
*       8 = U303/BB (-989 , -1033)
*       8 = U303/U211/VDD (-927.5 , -1089)
*       8 = U303/U210/VDD (-927.5 , -1038)
*       8 = U303/U215/VDD (-848.5 , -1085.5)
*       8 = U303/U213/VDD (-809 , -1037)
*       8 = U304/U211/VDD (-630 , -1089)
*       8 = U304/U210/VDD (-630 , -1038)
*       8 = U304/U215/VDD (-551 , -1085.5)
*       8 = U304/U213/VDD (-511.5 , -1037)
*       8 = U305/U211/VDD (-345.5 , -1089)
*       8 = U305/U210/VDD (-345.5 , -1038)
*       8 = U305/U215/VDD (-266.5 , -1085.5)
*       8 = U305/U213/VDD (-227 , -1037)
*       8 = U306/U210/VDD (-61 , -1038)
*       8 = U306/U211/VDD (-61 , -1089)
*       8 = U306/U215/VDD (18 , -1085.5)
*       8 = U306/U213/VDD (57.5 , -1037)
*       8 = U307/U215/VDD (302.5 , -1085.5)
*       8 = U307/U211/VDD (223.5 , -1089)
*       8 = U307/U210/VDD (223.5 , -1038)
*       8 = U307/U213/VDD (342 , -1037)
*       8 = U296/U211/VDD (507.5 , -1089)
*       8 = U296/U210/VDD (507.5 , -1038)
*       8 = U296/U215/VDD (586.5 , -1085.5)
*       8 = U296/U213/VDD (626 , -1037)
*       8 = U269/VDD (792 , -1038)
*       8 = U302/U234/VDD (-993 , -958.5)
*       8 = U302/U237/Vdd (-966 , -957.5)
*       8 = U302/U238/VDD (-871 , -961)
*       8 = U310/U211/VDD (-630 , -987)
*       8 = U310/U210/VDD (-630 , -936)
*       8 = U310/U215/VDD (-551 , -983.5)
*       8 = U310/U213/VDD (-511.5 , -935)
*       8 = U309/U228/VDD (-431.5 , -933.5)
*       8 = U309/U211/VDD (-345.5 , -987)
*       8 = U309/U210/VDD (-345.5 , -936)
*       8 = U309/U215/VDD (-266.5 , -983.5)
*       8 = U309/U213/VDD (-227 , -935)
*       8 = U308/U228/VDD (-147 , -933.5)
*       8 = U308/U210/VDD (-61 , -936)
*       8 = U308/U211/VDD (-61 , -987)
*       8 = U308/U215/VDD (18 , -983.5)
*       8 = U308/U213/VDD (57.5 , -935)
*       8 = U297/U228/VDD (137.5 , -933.5)
*       8 = U297/U215/VDD (302.5 , -983.5)
*       8 = U297/U211/VDD (223.5 , -987)
*       8 = U297/U210/VDD (223.5 , -936)
*       8 = U297/U213/VDD (342 , -935)
*       8 = U295/U228/VDD (421.5 , -933.5)
*       8 = U295/U210/VDD (507.5 , -936)
*       8 = U295/U211/VDD (507.5 , -987)
*       8 = U295/U215/VDD (586.5 , -983.5)
*       8 = U294/U228/VDD (706 , -933.5)
*       8 = U295/U213/VDD (626 , -935)
*       8 = U294/U210/VDD (792 , -936)
*       8 = U294/U211/VDD (792 , -987)
*       8 = U294/U215/VDD (871 , -983.5)
*       8 = U294/U213/VDD (910.5 , -935)
*       8 = U326/VddWell (-1685.5 , -862)
*       8 = U326/VddSel (-1684.5 , -862)
*       8 = U326/VddAct (-1682.5 , -862)
*       8 = U326/Vdd (-1617.5 , -862)
*       8 = U326/Vdd2 (-1682.5 , -862)
*       8 = U301/U234/VDD (-993 , -863.5)
*       8 = U301/U232/VDD (-906.9 , -865.9)
*       8 = U242/U229/VDD (-730.5 , -836.5)
*       8 = U242/U228/VDD (-716 , -888.5)
*       8 = U242/U211/VDD (-620.5 , -891)
*       8 = U242/U210/VDD (-620.5 , -840)
*       8 = U242/U215/VDD (-541.5 , -887.5)
*       8 = U242/U213/VDD (-502 , -839)
*       8 = U244/U229/VDD (-446 , -836.5)
*       8 = U244/U228/VDD (-431.5 , -888.5)
*       8 = U244/U211/VDD (-336 , -891)
*       8 = U244/U210/VDD (-336 , -840)
*       8 = U244/U215/VDD (-257 , -887.5)
*       8 = U244/U213/VDD (-217.5 , -839)
*       8 = U246/U229/VDD (-161.5 , -836.5)
*       8 = U246/U228/VDD (-147 , -888.5)
*       8 = U246/U211/VDD (-51.5 , -891)
*       8 = U246/U210/VDD (-51.5 , -840)
*       8 = U246/U215/VDD (27.5 , -887.5)
*       8 = U246/U213/VDD (67 , -839)
*       8 = U248/U229/VDD (123 , -836.5)
*       8 = U248/U228/VDD (137.5 , -888.5)
*       8 = U248/U211/VDD (233 , -891)
*       8 = U248/U210/VDD (233 , -840)
*       8 = U250/U229/VDD (407 , -836.5)
*       8 = U248/U213/VDD (351.5 , -839)
*       8 = U248/U215/VDD (312 , -887.5)
*       8 = U250/U228/VDD (421.5 , -888.5)
*       8 = U250/U215/VDD (596 , -887.5)
*       8 = U250/U211/VDD (517 , -891)
*       8 = U250/U210/VDD (517 , -840)
*       8 = U252/U229/VDD (691.5 , -836.5)
*       8 = U250/U213/VDD (635.5 , -839)
*       8 = U252/U228/VDD (706 , -888.5)
*       8 = U252/U210/VDD (801.5 , -840)
*       8 = U252/U211/VDD (801.5 , -891)
*       8 = U252/U215/VDD (880.5 , -887.5)
*       8 = U252/U213/VDD (920 , -839)
*       8 = U342/VddWell (1491.5 , -866)
*       8 = U342/VddSel (1492.5 , -866)
*       8 = U342/VddAct (1494.5 , -866)
*       8 = U342/Vdd (1494.5 , -866)
*       8 = U342/Vdd2 (1559.5 , -866)
*       8 = U300/U234/VDD (-993 , -767.5)
*       8 = U300/U232/VDD (-906.9 , -769.9)
*       8 = U241/U229/VDD (-730.5 , -740.5)
*       8 = U241/U228/VDD (-716 , -792.5)
*       8 = U241/U211/VDD (-620.5 , -795)
*       8 = U241/U210/VDD (-620.5 , -744)
*       8 = U241/U215/VDD (-541.5 , -791.5)
*       8 = U241/U213/VDD (-502 , -743)
*       8 = U243/U229/VDD (-446 , -740.5)
*       8 = U243/U228/VDD (-431.5 , -792.5)
*       8 = U243/U211/VDD (-336 , -795)
*       8 = U243/U210/VDD (-336 , -744)
*       8 = U243/U215/VDD (-257 , -791.5)
*       8 = U243/U213/VDD (-217.5 , -743)
*       8 = U245/U229/VDD (-161.5 , -740.5)
*       8 = U245/U228/VDD (-147 , -792.5)
*       8 = U245/U211/VDD (-51.5 , -795)
*       8 = U245/U210/VDD (-51.5 , -744)
*       8 = U245/U215/VDD (27.5 , -791.5)
*       8 = U245/U213/VDD (67 , -743)
*       8 = U247/U229/VDD (123 , -740.5)
*       8 = U247/U228/VDD (137.5 , -792.5)
*       8 = U247/U211/VDD (233 , -795)
*       8 = U247/U210/VDD (233 , -744)
*       8 = U249/U229/VDD (407 , -740.5)
*       8 = U247/U213/VDD (351.5 , -743)
*       8 = U247/U215/VDD (312 , -791.5)
*       8 = U249/U228/VDD (421.5 , -792.5)
*       8 = U249/U215/VDD (596 , -791.5)
*       8 = U249/U211/VDD (517 , -795)
*       8 = U249/U210/VDD (517 , -744)
*       8 = U251/U229/VDD (691.5 , -740.5)
*       8 = U249/U213/VDD (635.5 , -743)
*       8 = U251/U228/VDD (706 , -792.5)
*       8 = U251/U210/VDD (801.5 , -744)
*       8 = U251/U211/VDD (801.5 , -795)
*       8 = U251/U215/VDD (880.5 , -791.5)
*       8 = U251/U213/VDD (920 , -743)
*       8 = U299/U234/VDD (-993 , -672.5)
*       8 = U299/U232/VDD (-906.9 , -674.9)
*       8 = U281/U237/Vdd (-689 , -671.5)
*       8 = U281/U234/VDD (-716 , -672.5)
*       8 = U281/U238/VDD (-594 , -675)
*       8 = U279/U229/VDD (-446 , -644.5)
*       8 = U279/U228/VDD (-431.5 , -696.5)
*       8 = U279/U211/VDD (-336 , -699)
*       8 = U279/U210/VDD (-336 , -648)
*       8 = U279/U213/VDD (-217.5 , -647)
*       8 = U279/U215/VDD (-257 , -695.5)
*       8 = U282/U237/Vdd (-107.5 , -670.5)
*       8 = U282/U234/VDD (-134.5 , -671.5)
*       8 = U282/U238/VDD (-12.5 , -674)
*       8 = U283/U237/Vdd (177 , -670.5)
*       8 = U283/U234/VDD (150 , -671.5)
*       8 = U283/U238/VDD (272 , -674)
*       8 = U284/U237/Vdd (461 , -670.5)
*       8 = U284/U234/VDD (434 , -671.5)
*       8 = U284/U238/VDD (556 , -674)
*       8 = U285/U237/Vdd (745.5 , -670.5)
*       8 = U285/U234/VDD (718.5 , -671.5)
*       8 = U285/U238/VDD (840.5 , -674)
*       8 = U298/U234/VDD (-993 , -594.5)
*       8 = U298/U232/VDD (-906.9 , -596.9)
*       8 = U298/U232/A (-874.9 , -598.4)
*       8 = U298/AA (-875 , -593.5)
*       8 = U287/U240/VDD (-728 , -593.5)
*       8 = U287/U239/VDD (-753 , -594.5)
*       8 = U293/U237/Vdd (-404.5 , -592.5)
*       8 = U293/U234/VDD (-431.5 , -593.5)
*       8 = U293/U238/VDD (-309.5 , -596)
*       8 = U293/U238/A (-277.5 , -597.5)
*       8 = U293/AA (-277.5 , -593.5)
*       8 = U288/U240/VDD (-146.5 , -592.5)
*       8 = U288/U239/VDD (-171.5 , -593.5)
*       8 = U289/U240/VDD (138 , -592.5)
*       8 = U289/U239/VDD (113 , -593.5)
*       8 = U290/U239/VDD (397 , -593.5)
*       8 = U290/U240/VDD (422 , -592.5)
*       8 = U291/U240/VDD (706.5 , -592.5)
*       8 = U291/U239/VDD (681.5 , -593.5)
*       8 = U327/VddWell (-1685.5 , -426)
*       8 = U327/VddSel (-1684.5 , -426)
*       8 = U327/VddAct (-1682.5 , -426)
*       8 = U327/Vdd (-1617.5 , -426)
*       8 = U327/Vdd2 (-1682.5 , -426)
*       8 = U343/VddWell (1491.5 , -430)
*       8 = U343/VddSel (1492.5 , -430)
*       8 = U343/VddAct (1494.5 , -430)
*       8 = U343/Vdd (1494.5 , -430)
*       8 = U343/Vdd2 (1559.5 , -430)
*       8 = U328/VddWell (-1685.5 , 10)
*       8 = U328/VddSel (-1684.5 , 10)
*       8 = U328/VddAct (-1682.5 , 10)
*       8 = U328/Vdd (-1617.5 , 10)
*       8 = U328/Vdd2 (-1682.5 , 10)
*       8 = U329/VddWell (1491.5 , 10)
*       8 = U329/VddSel (1492.5 , 10)
*       8 = U329/VddAct (1494.5 , 10)
*       8 = U329/Vdd (1494.5 , 10)
*       8 = U329/Vdd2 (1559.5 , 10)
*       8 = U322/VddWell (-1685.5 , 446)
*       8 = U322/VddSel (-1684.5 , 446)
*       8 = U322/VddAct (-1682.5 , 446)
*       8 = U322/Vdd (-1617.5 , 446)
*       8 = U322/Vdd2 (-1682.5 , 446)
*       8 = U313/VddWell (-1557.5 , 443)
*       8 = U313/VddSel (-1557.5 , 444)
*       8 = U313/VddAct (-1557.5 , 446)
*       8 = U313/Vdd (-1557.5 , 446)
*       8 = U315/VddWell (-1121.5 , 443)
*       8 = U315/VddSel (-1121.5 , 444)
*       8 = U315/VddAct (-1121.5 , 446)
*       8 = U315/Vdd (-1121.5 , 446)
*       8 = U316/VddWell (-685.5 , 443)
*       8 = U316/VddSel (-685.5 , 444)
*       8 = U316/VddAct (-685.5 , 446)
*       8 = U316/Vdd (-685.5 , 446)
*       8 = U317/VddWell (-249.5 , 443)
*       8 = U317/VddSel (-249.5 , 444)
*       8 = U317/VddAct (-249.5 , 446)
*       8 = U317/Vdd (-249.5 , 446)
*       8 = U318/VddWell (186.5 , 443)
*       8 = U318/VddSel (186.5 , 444)
*       8 = U318/VddAct (186.5 , 446)
*       8 = U318/Vdd (186.5 , 446)
*       8 = U319/VddWell (622.5 , 443)
*       8 = U319/VddSel (622.5 , 444)
*       8 = U319/VddAct (622.5 , 446)
*       8 = U319/Vdd (622.5 , 446)
*       8 = U320/VddWell (1058.5 , 443)
*       8 = U320/VddSel (1058.5 , 444)
*       8 = U320/VddAct (1058.5 , 446)
*       8 = U320/Vdd (1058.5 , 446)
*       8 = U323/VddWell (1491.5 , 446)
*       8 = U323/VddSel (1492.5 , 446)
*       8 = U323/VddAct (1494.5 , 446)
*       8 = U323/Vdd (1494.5 , 446)
*       8 = U323/Vdd2 (1559.5 , 446)
*       8 = U313/Vdd2 (-1557.5 , 511)
*       8 = U315/Vdd2 (-1121.5 , 511)
*       8 = U316/Vdd2 (-685.5 , 511)
*       8 = U317/Vdd2 (-249.5 , 511)
*       8 = U318/Vdd2 (186.5 , 511)
*       8 = U319/Vdd2 (622.5 , 511)
*       8 = U320/Vdd2 (1058.5 , 511)
*       12 = U329/Gnd (1494.5 , 88)
*       12 = U310/U211/GND (-639 , -1017.5)
*       12 = U303/U210/GND (-936.5 , -1068.5)
*       12 = U303/U211/GND (-936.5 , -1119.5)
*       12 = U331/GndSel (-1557.5 , -2432)
*       12 = U331/GndAct (-1557.5 , -2430)
*       12 = U330/GndSel (-1557.5 , -2432)
*       12 = U330/GndAct (-1557.5 , -2430)
*       12 = U331/Gnd2 (-1557.5 , -2430)
*       12 = U330/Gnd2 (-1557.5 , -2430)
*       12 = U332/GndSel (-1121.5 , -2432)
*       12 = U332/GndAct (-1121.5 , -2430)
*       12 = U332/Gnd2 (-1121.5 , -2430)
*       12 = U333/GndSel (-685.5 , -2432)
*       12 = U333/GndAct (-685.5 , -2430)
*       12 = U333/Gnd2 (-685.5 , -2430)
*       12 = U334/GndSel (-249.5 , -2432)
*       12 = U334/GndAct (-249.5 , -2430)
*       12 = U334/Gnd2 (-249.5 , -2430)
*       12 = U335/GndSel (186.5 , -2432)
*       12 = U335/GndAct (186.5 , -2430)
*       12 = U335/Gnd2 (186.5 , -2430)
*       12 = U336/GndSel (622.5 , -2432)
*       12 = U336/GndAct (622.5 , -2430)
*       12 = U336/Gnd2 (622.5 , -2430)
*       12 = U337/GndSel (1058.5 , -2432)
*       12 = U337/GndAct (1058.5 , -2430)
*       12 = U337/Gnd2 (1058.5 , -2430)
*       12 = U338/GndSel (1494.5 , -2432)
*       12 = U338/GndAct (1494.5 , -2430)
*       12 = U338/Gnd2 (1494.5 , -2430)
*       12 = U331/Gnd (-1557.5 , -2365)
*       12 = U330/Gnd (-1557.5 , -2365)
*       12 = U332/Gnd (-1121.5 , -2365)
*       12 = U333/Gnd (-685.5 , -2365)
*       12 = U334/Gnd (-249.5 , -2365)
*       12 = U335/Gnd (186.5 , -2365)
*       12 = U336/Gnd (622.5 , -2365)
*       12 = U337/Gnd (1058.5 , -2365)
*       12 = U338/Gnd (1494.5 , -2365)
*       12 = U344/GndSel (-1815.5 , -2170)
*       12 = U344/GndAct (-1813.5 , -2170)
*       12 = U344/Gnd2 (-1813.5 , -2170)
*       12 = U344/Gnd (-1748.5 , -2170)
*       12 = U339/GndSel (1623.5 , -2174)
*       12 = U339/GndAct (1625.5 , -2174)
*       12 = U339/Gnd (1625.5 , -2174)
*       12 = U339/Gnd2 (1690.5 , -2174)
*       12 = U324/GndSel (-1815.5 , -1734)
*       12 = U324/GndAct (-1813.5 , -1734)
*       12 = U324/Gnd2 (-1813.5 , -1734)
*       12 = U324/Gnd (-1748.5 , -1734)
*       12 = U340/GndSel (1623.5 , -1738)
*       12 = U340/GndAct (1625.5 , -1738)
*       12 = U340/Gnd (1625.5 , -1738)
*       12 = U340/Gnd2 (1690.5 , -1738)
*       12 = U325/GndSel (-1815.5 , -1298)
*       12 = U325/GndAct (-1813.5 , -1298)
*       12 = U325/Gnd2 (-1813.5 , -1298)
*       12 = U325/Gnd (-1748.5 , -1298)
*       12 = U341/GndSel (1623.5 , -1302)
*       12 = U341/GndAct (1625.5 , -1302)
*       12 = U341/Gnd (1625.5 , -1302)
*       12 = U341/Gnd2 (1690.5 , -1302)
*       12 = U303/U215/GND (-834.5 , -1120.5)
*       12 = U304/U211/GND (-639 , -1119.5)
*       12 = U304/U215/GND (-537 , -1120.5)
*       12 = U305/U211/GND (-354.5 , -1119.5)
*       12 = U305/U215/GND (-252.5 , -1120.5)
*       12 = U306/U211/GND (-70 , -1119.5)
*       12 = U306/U215/GND (32 , -1120.5)
*       12 = U307/U211/GND (214.5 , -1119.5)
*       12 = U307/U215/GND (316.5 , -1120.5)
*       12 = U296/U211/GND (498.5 , -1119.5)
*       12 = U296/U215/GND (600.5 , -1120.5)
*       12 = U303/U213/GND (-817.5 , -1069)
*       12 = U304/U210/GND (-639 , -1068.5)
*       12 = U304/U213/GND (-520 , -1069)
*       12 = U310/U215/GND (-537 , -1018.5)
*       12 = U309/U211/GND (-354.5 , -1017.5)
*       12 = U305/U210/GND (-354.5 , -1068.5)
*       12 = U305/U213/GND (-235.5 , -1069)
*       12 = U309/U215/GND (-252.5 , -1018.5)
*       12 = U306/U210/GND (-70 , -1068.5)
*       12 = U308/U211/GND (-70 , -1017.5)
*       12 = U306/U213/GND (49 , -1069)
*       12 = U308/U215/GND (32 , -1018.5)
*       12 = U297/U211/GND (214.5 , -1017.5)
*       12 = U307/U210/GND (214.5 , -1068.5)
*       12 = U307/U213/GND (333.5 , -1069)
*       12 = U297/U215/GND (316.5 , -1018.5)
*       12 = U296/U210/GND (498.5 , -1068.5)
*       12 = U295/U211/GND (498.5 , -1017.5)
*       12 = U295/U215/GND (600.5 , -1018.5)
*       12 = U296/U213/GND (617.5 , -1069)
*       12 = U294/U211/GND (783 , -1017.5)
*       12 = U269/GND (783 , -1068.5)
*       12 = U294/U215/GND (885 , -1018.5)
*       12 = U302/U234/GND (-1042.5 , -993)
*       12 = U302/U237/GND (-967.5 , -992)
*       12 = U302/U238/GND (-880 , -991.5)
*       12 = U242/U228/GND (-765.5 , -923)
*       12 = U310/U228/GND (-765.5 , -968)
*       12 = U310/U210/GND (-639 , -966.5)
*       12 = U242/U211/GND (-629.5 , -921.5)
*       12 = U242/U215/GND (-527.5 , -922.5)
*       12 = U310/U213/GND (-520 , -967)
*       12 = U244/U228/GND (-481 , -923)
*       12 = U309/U228/GND (-481 , -968)
*       12 = U309/U210/GND (-354.5 , -966.5)
*       12 = U244/U211/GND (-345 , -921.5)
*       12 = U246/U228/GND (-196.5 , -923)
*       12 = U244/U215/GND (-243 , -922.5)
*       12 = U309/U213/GND (-235.5 , -967)
*       12 = U308/U228/GND (-196.5 , -968)
*       12 = U308/U210/GND (-70 , -966.5)
*       12 = U246/U211/GND (-60.5 , -921.5)
*       12 = U248/U228/GND (88 , -923)
*       12 = U246/U215/GND (41.5 , -922.5)
*       12 = U308/U213/GND (49 , -967)
*       12 = U297/U228/GND (88 , -968)
*       12 = U248/U211/GND (224 , -921.5)
*       12 = U297/U210/GND (214.5 , -966.5)
*       12 = U297/U213/GND (333.5 , -967)
*       12 = U295/U228/GND (372 , -968)
*       12 = U250/U228/GND (372 , -923)
*       12 = U248/U215/GND (326 , -922.5)
*       12 = U250/U211/GND (508 , -921.5)
*       12 = U295/U210/GND (498.5 , -966.5)
*       12 = U250/U215/GND (610 , -922.5)
*       12 = U252/U228/GND (656.5 , -923)
*       12 = U294/U228/GND (656.5 , -968)
*       12 = U295/U213/GND (617.5 , -967)
*       12 = U294/U210/GND (783 , -966.5)
*       12 = U252/U211/GND (792.5 , -921.5)
*       12 = U252/U215/GND (894.5 , -922.5)
*       12 = U294/U213/GND (902 , -967)
*       12 = U326/GndSel (-1815.5 , -862)
*       12 = U326/GndAct (-1813.5 , -862)
*       12 = U326/Gnd2 (-1813.5 , -862)
*       12 = U326/Gnd (-1748.5 , -862)
*       12 = U301/U234/GND (-1042.5 , -898)
*       12 = U301/U232/GND (-915.9 , -896.4)
*       12 = U241/U228/GND (-765.5 , -827)
*       12 = U242/U229/GND (-716.5 , -871.5)
*       12 = U242/U210/GND (-629.5 , -870.5)
*       12 = U241/U211/GND (-629.5 , -825.5)
*       12 = U241/U215/GND (-527.5 , -826.5)
*       12 = U242/U213/GND (-510.5 , -871)
*       12 = U243/U228/GND (-481 , -827)
*       12 = U244/U229/GND (-432 , -871.5)
*       12 = U244/U210/GND (-345 , -870.5)
*       12 = U243/U211/GND (-345 , -825.5)
*       12 = U245/U228/GND (-196.5 , -827)
*       12 = U243/U215/GND (-243 , -826.5)
*       12 = U244/U213/GND (-226 , -871)
*       12 = U246/U229/GND (-147.5 , -871.5)
*       12 = U246/U210/GND (-60.5 , -870.5)
*       12 = U245/U211/GND (-60.5 , -825.5)
*       12 = U247/U228/GND (88 , -827)
*       12 = U245/U215/GND (41.5 , -826.5)
*       12 = U246/U213/GND (58.5 , -871)
*       12 = U248/U229/GND (137 , -871.5)
*       12 = U247/U211/GND (224 , -825.5)
*       12 = U248/U210/GND (224 , -870.5)
*       12 = U249/U228/GND (372 , -827)
*       12 = U247/U215/GND (326 , -826.5)
*       12 = U248/U213/GND (343 , -871)
*       12 = U249/U211/GND (508 , -825.5)
*       12 = U250/U229/GND (421 , -871.5)
*       12 = U250/U210/GND (508 , -870.5)
*       12 = U249/U215/GND (610 , -826.5)
*       12 = U252/U229/GND (705.5 , -871.5)
*       12 = U250/U213/GND (627 , -871)
*       12 = U251/U228/GND (656.5 , -827)
*       12 = U252/U210/GND (792.5 , -870.5)
*       12 = U251/U211/GND (792.5 , -825.5)
*       12 = U251/U215/GND (894.5 , -826.5)
*       12 = U252/U213/GND (911.5 , -871)
*       12 = U342/GndSel (1623.5 , -866)
*       12 = U342/GndAct (1625.5 , -866)
*       12 = U342/Gnd (1625.5 , -866)
*       12 = U342/Gnd2 (1690.5 , -866)
*       12 = U299/U234/GND (-1042.5 , -707)
*       12 = U300/U234/GND (-1042.5 , -802)
*       12 = U300/U232/GND (-915.9 , -800.4)
*       12 = U299/U232/GND (-915.9 , -705.4)
*       12 = U241/U229/GND (-716.5 , -775.5)
*       12 = U281/U237/GND (-690.5 , -706)
*       12 = U281/U234/GND (-765.5 , -707)
*       12 = U281/U238/GND (-603 , -705.5)
*       12 = U241/U210/GND (-629.5 , -774.5)
*       12 = U241/U213/GND (-510.5 , -775)
*       12 = U243/U229/GND (-432 , -775.5)
*       12 = U279/U228/GND (-481 , -731)
*       12 = U279/U211/GND (-345 , -729.5)
*       12 = U243/U210/GND (-345 , -774.5)
*       12 = U243/U213/GND (-226 , -775)
*       12 = U279/U215/GND (-243 , -730.5)
*       12 = U282/U234/GND (-184 , -706)
*       12 = U245/U229/GND (-147.5 , -775.5)
*       12 = U245/U210/GND (-60.5 , -774.5)
*       12 = U283/U234/GND (100.5 , -706)
*       12 = U245/U213/GND (58.5 , -775)
*       12 = U247/U229/GND (137 , -775.5)
*       12 = U247/U210/GND (224 , -774.5)
*       12 = U284/U234/GND (384.5 , -706)
*       12 = U247/U213/GND (343 , -775)
*       12 = U249/U229/GND (421 , -775.5)
*       12 = U249/U210/GND (508 , -774.5)
*       12 = U285/U234/GND (669 , -706)
*       12 = U251/U229/GND (705.5 , -775.5)
*       12 = U249/U213/GND (627 , -775)
*       12 = U251/U210/GND (792.5 , -774.5)
*       12 = U251/U213/GND (911.5 , -775)
*       12 = U298/U234/GND (-1042.5 , -629)
*       12 = U298/U232/GND (-915.9 , -627.4)
*       12 = U287/U240/GND (-714 , -628.5)
*       12 = U287/U239/GND (-723.5 , -628.5)
*       12 = U279/U229/GND (-432 , -679.5)
*       12 = U293/U237/GND (-406 , -627)
*       12 = U293/U234/GND (-481 , -628)
*       12 = U293/U238/GND (-318.5 , -626.5)
*       12 = U279/U210/GND (-345 , -678.5)
*       12 = U279/U213/GND (-226 , -679)
*       12 = U282/U237/GND (-109 , -705)
*       12 = U288/U240/GND (-132.5 , -627.5)
*       12 = U288/U239/GND (-142 , -627.5)
*       12 = U282/U238/GND (-21.5 , -704.5)
*       12 = U283/U237/GND (175.5 , -705)
*       12 = U289/U240/GND (152 , -627.5)
*       12 = U289/U239/GND (142.5 , -627.5)
*       12 = U283/U238/GND (263 , -704.5)
*       12 = U284/U237/GND (459.5 , -705)
*       12 = U290/U240/GND (436 , -627.5)
*       12 = U290/U239/GND (426.5 , -627.5)
*       12 = U284/U238/GND (547 , -704.5)
*       12 = U291/U239/GND (711 , -627.5)
*       12 = U285/U237/GND (744 , -705)
*       12 = U291/U240/GND (720.5 , -627.5)
*       12 = U285/U238/GND (831.5 , -704.5)
*       12 = U327/GndSel (-1815.5 , -426)
*       12 = U327/GndAct (-1813.5 , -426)
*       12 = U327/Gnd2 (-1813.5 , -426)
*       12 = U327/Gnd (-1748.5 , -426)
*       12 = U343/GndSel (1623.5 , -430)
*       12 = U343/GndAct (1625.5 , -430)
*       12 = U343/Gnd (1625.5 , -430)
*       12 = U343/Gnd2 (1690.5 , -430)
*       12 = U328/GndSel (-1815.5 , 10)
*       12 = U328/GndAct (-1813.5 , 10)
*       12 = U328/Gnd2 (-1813.5 , 10)
*       12 = U328/Gnd (-1748.5 , 10)
*       12 = U329/GndSel (1623.5 , 10)
*       12 = U329/GndAct (1625.5 , 10)
*       12 = U329/Gnd2 (1690.5 , 10)
*       12 = U322/GndSel (-1815.5 , 446)
*       12 = U322/GndAct (-1813.5 , 446)
*       12 = U322/Gnd2 (-1813.5 , 446)
*       12 = U322/Gnd (-1748.5 , 446)
*       12 = U323/GndSel (1623.5 , 446)
*       12 = U323/GndAct (1625.5 , 446)
*       12 = U323/Gnd (1625.5 , 446)
*       12 = U323/Gnd2 (1690.5 , 446)
*       12 = U313/GndSel (-1557.5 , 575)
*       12 = U313/GndAct (-1557.5 , 577)
*       12 = U313/Gnd (-1557.5 , 577)
*       12 = U315/GndSel (-1121.5 , 575)
*       12 = U315/GndAct (-1121.5 , 577)
*       12 = U315/Gnd (-1121.5 , 577)
*       12 = U316/GndSel (-685.5 , 575)
*       12 = U316/GndAct (-685.5 , 577)
*       12 = U316/Gnd (-685.5 , 577)
*       12 = U317/GndSel (-249.5 , 575)
*       12 = U317/GndAct (-249.5 , 577)
*       12 = U317/Gnd (-249.5 , 577)
*       12 = U318/GndSel (186.5 , 575)
*       12 = U318/GndAct (186.5 , 577)
*       12 = U318/Gnd (186.5 , 577)
*       12 = U319/GndSel (622.5 , 575)
*       12 = U319/GndAct (622.5 , 577)
*       12 = U319/Gnd (622.5 , 577)
*       12 = U320/GndSel (1058.5 , 575)
*       12 = U320/GndAct (1058.5 , 577)
*       12 = U320/Gnd (1058.5 , 577)
*       12 = U313/Gnd2 (-1557.5 , 642)
*       12 = U315/Gnd2 (-1121.5 , 642)
*       12 = U316/Gnd2 (-685.5 , 642)
*       12 = U317/Gnd2 (-249.5 , 642)
*       12 = U318/Gnd2 (186.5 , 642)
*       12 = U319/Gnd2 (622.5 , 642)
*       12 = U320/Gnd2 (1058.5 , 642)
*       17 = U318/DataInB (333.5 , 446)
*       18 = U297/U228/INPUTB (119 , -962)
*       18 = U248/U228/INPUTB (119 , -917)
*       18 = U248/Y (120.5 , -836.5)
*       18 = U247/U228/INPUTB (119 , -821)
*       18 = U247/Y (120.5 , -740.5)
*       18 = U289/U239/B (134 , -615)
*       18 = U283/U234/INPUTB (131.5 , -700)
*       18 = U283/Y (133.5 , -671)
*       18 = U289/Y (133.5 , -591)
*       18 = Y2 (133.5 , -591)
*       18 = U318/DataIn (309.5 , 446)
*       24 = U316/DataInB (-538.5 , 446)
*       31 = U320/DataInB (1205.5 , 446)
*       33 = U319/DataInB (769.5 , 446)
*       35 = U317/DataInB (-102.5 , 446)
*       37 = U309/U228/INPUTB (-450 , -962)
*       37 = U244/U228/INPUTB (-450 , -917)
*       37 = U244/Y (-448.5 , -836.5)
*       37 = U243/U228/INPUTB (-450 , -821)
*       37 = U279/U228/INPUTB (-450 , -725)
*       37 = U243/Y (-448.5 , -740.5)
*       37 = U293/U234/INPUTB (-450 , -622)
*       37 = U279/Y (-448.5 , -644.5)
*       37 = U293/Y (-448 , -593)
*       37 = Y4 (-448 , -591)
*       37 = U316/DataIn (-562.5 , 446)
*       38 = U315/DataInB (-974.5 , 446)
*       39 = U313/DataInB (-1410.5 , 446)
*       40 = U310/U228/INPUTB (-734.5 , -962)
*       40 = U242/U228/INPUTB (-734.5 , -917)
*       40 = U242/Y (-733 , -836.5)
*       40 = U241/U228/INPUTB (-734.5 , -821)
*       40 = U241/Y (-733 , -740.5)
*       40 = U287/U239/B (-732 , -616)
*       40 = U281/U234/INPUTB (-734.5 , -701)
*       40 = U281/Y (-732.5 , -672)
*       40 = U287/Y (-732.5 , -592)
*       40 = Y5 (-732.5 , -592)
*       40 = U315/DataIn (-998.5 , 446)
*       41 = U302/U234/INPUTB (-1011.5 , -987)
*       41 = U302/Y (-1009.5 , -958)
*       41 = U301/U234/INPUTB (-1011.5 , -892)
*       41 = U301/Y (-1009.5 , -863)
*       41 = U300/U234/INPUTB (-1011.5 , -796)
*       41 = U300/Y (-1009.5 , -767)
*       41 = U299/U234/INPUTB (-1011.5 , -701)
*       41 = U299/Y (-1009.5 , -672)
*       41 = U298/U234/INPUTB (-1011.5 , -623)
*       41 = U298/Y (-1009.5 , -594)
*       41 = Y6 (-1009.5 , -592)
*       41 = U313/DataIn (-1434.5 , 446)
*       45 = U328/DataIn (-1557.5 , 133)
*       45 = U298/U234/INPUTA (-1067 , -625)
*       45 = U298/X (-1072 , -611)
*       45 = X0 (-1072.5 , -613)
*       45 = U287/U239/A (-758.5 , -616)
*       45 = U287/X (-764.5 , -611)
*       45 = U293/U234/INPUTA (-505.5 , -624)
*       45 = U293/X (-510.5 , -610.5)
*       45 = U288/U239/A (-177 , -615)
*       45 = U288/X (-183 , -610)
*       45 = U289/U239/A (107.5 , -615)
*       45 = U289/X (101.5 , -610)
*       45 = U290/U239/A (391.5 , -615)
*       45 = U290/X (385.5 , -610)
*       45 = U291/U239/A (676 , -615)
*       45 = U291/X (670 , -610)
*       46 = U328/DataInB (-1557.5 , 157)
*       47 = U328/DataInUnBuf (-1557.5 , 173)
*       54 = U327/DataIn (-1557.5 , -303)
*       54 = U299/U234/INPUTA (-1067 , -703)
*       54 = U299/X (-1072 , -689)
*       54 = X1 (-1073 , -691.5)
*       54 = U281/U234/INPUTA (-790 , -703)
*       54 = U281/X (-795 , -689.5)
*       54 = U279/U228/INPUTA (-505.5 , -727)
*       54 = U279/X (-510.5 , -688)
*       54 = U282/U234/INPUTA (-208.5 , -702)
*       54 = U282/X (-213.5 , -688.5)
*       54 = U283/U234/INPUTA (76 , -702)
*       54 = U283/X (71 , -688.5)
*       54 = U284/U234/INPUTA (360 , -702)
*       54 = U284/X (355 , -688.5)
*       54 = U285/U234/INPUTA (644.5 , -702)
*       54 = U285/X (639.5 , -688.5)
*       58 = U327/DataInB (-1557.5 , -279)
*       59 = U327/DataInUnBuf (-1557.5 , -263)
*       62 = U293/U237/vout (-385.5 , -616)
*       62 = U293/U238/B (-371 , -599.5)
*       70 = U291/U239/OUT (689.5 , -626.5)
*       70 = U291/U240/vin (728 , -614.5)
*       71 = U285/U237/vin (736 , -693)
*       71 = U285/U234/OUTPUT (725 , -684.5)
*       72 = U291/U240/vout (713.5 , -613)
*       72 = P0 (915.5 , -656)
*       72 = U343/DataOut (1494.5 , -169)
*       73 = U294/U228/INPUTB (687.5 , -962)
*       73 = U252/U228/INPUTB (687.5 , -917)
*       73 = U252/Y (689 , -836.5)
*       73 = U251/U228/INPUTB (687.5 , -821)
*       73 = U251/Y (689 , -740.5)
*       73 = U291/U239/B (702.5 , -615)
*       73 = U285/U234/INPUTB (700 , -700)
*       73 = U285/Y (702 , -671)
*       73 = U291/Y (702 , -591)
*       73 = Y0 (702 , -591)
*       73 = U320/DataIn (1181.5 , 446)
*       82 = U290/U240/vout (429 , -613)
*       82 = U285/U238/A (872.5 , -675.5)
*       82 = U285/AA (872.5 , -671.5)
*       83 = U295/U228/INPUTB (403 , -962)
*       83 = U250/U228/INPUTB (403 , -917)
*       83 = U250/Y (404.5 , -836.5)
*       83 = U249/U228/INPUTB (403 , -821)
*       83 = U249/Y (404.5 , -740.5)
*       83 = U290/U239/B (418 , -615)
*       83 = U284/U234/INPUTB (415.5 , -700)
*       83 = U284/Y (417.5 , -671)
*       83 = U290/Y (417.5 , -591)
*       83 = Y1 (417.5 , -591)
*       83 = U319/DataIn (745.5 , 446)
*       84 = U290/U239/OUT (405 , -626.5)
*       84 = U290/U240/vin (443.5 , -614.5)
*       85 = U284/U237/vin (451.5 , -693)
*       85 = U284/U234/OUTPUT (440.5 , -684.5)
*       91 = U289/U239/OUT (121 , -626.5)
*       91 = U289/U240/vin (159.5 , -614.5)
*       94 = U289/U240/vout (145 , -613)
*       94 = U284/U238/A (588 , -675.5)
*       94 = U284/AA (588 , -671.5)
*       95 = U283/U237/vin (167.5 , -693)
*       95 = U283/U234/OUTPUT (156.5 , -684.5)
*       101 = U288/U239/OUT (-163.5 , -626.5)
*       101 = U288/U240/vin (-125 , -614.5)
*       104 = U288/U240/vout (-139.5 , -613)
*       104 = U283/U238/A (304 , -675.5)
*       104 = U283/AA (304 , -671.5)
*       105 = U282/U237/vin (-117 , -693)
*       105 = U282/U234/OUTPUT (-128 , -684.5)
*       108 = U279/U210/A (-304 , -649.5)
*       108 = U279/AA (-304 , -643.5)
*       108 = U293/Carry (-263 , -629.5)
*       108 = U293/U238/C (-263 , -597)
*       114 = U279/U210/C (-289.5 , -649)
*       114 = U279/U213/A (-253 , -651)
*       116 = U293/Sum (-379 , -630)
*       116 = U282/U238/A (19.5 , -675.5)
*       116 = U282/AA (19.5 , -671.5)
*       116 = U293/U238/S (-379 , -599)
*       120 = U279/U210/B (-397.5 , -651.5)
*       120 = U279/BB (-397.5 , -643)
*       120 = U279/U229/vout (-439 , -665)
*       121 = U293/U234/OUTPUT (-425 , -606.5)
*       121 = U293/U237/vin (-414 , -615)
*       128 = U287/U239/OUT (-745 , -627.5)
*       128 = U287/U240/vin (-706.5 , -615.5)
*       130 = U281/U237/vout (-670 , -695)
*       130 = U281/U238/B (-655.5 , -678.5)
*       132 = U287/U240/vout (-721 , -614)
*       132 = U279/U211/A (-304 , -700.5)
*       132 = U279/CC (-378.5 , -643)
*       143 = U298/Sum (-976.5 , -630)
*       143 = U281/U238/A (-562 , -676.5)
*       143 = U281/AA (-562 , -672.5)
*       143 = U298/U232/S (-976.4 , -599.9)
*       144 = U299/U232/B (-968.4 , -678.4)
*       144 = U299/U234/OUTPUT (-986.5 , -685.5)
*       146 = U298/U234/OUTPUT (-986.5 , -607.5)
*       146 = U298/U232/B (-968.4 , -600.4)
*       153 = U251/U213/A (884.5 , -747)
*       153 = U251/U210/C (848 , -745)
*       160 = U285/Sum (771 , -708)
*       160 = P1 (915.5 , -715)
*       160 = U285/U238/S (771 , -677)
*       160 = U342/DataOut (1494.5 , -605)
*       161 = U285/U237/vout (764.5 , -694)
*       161 = U285/U238/B (779 , -677.5)
*       163 = U285/Carry (887 , -707.5)
*       163 = U251/U210/A (833.5 , -745.5)
*       163 = U251/AA (833.5 , -739.5)
*       163 = U285/U238/C (887 , -675)
*       164 = U251/U229/vout (698.5 , -761)
*       164 = U251/U210/B (740 , -747.5)
*       164 = U251/BB (740 , -739)
*       165 = U251/U228/OUTPUT (712.5 , -805.5)
*       165 = U251/U229/vin (713 , -762.5)
*       167 = U249/U213/A (600 , -747)
*       167 = U249/U210/C (563.5 , -745)
*       172 = U284/Sum (486.5 , -708)
*       172 = U251/CC (759 , -739)
*       172 = U251/U211/A (833.5 , -796.5)
*       172 = U284/U238/S (486.5 , -677)
*       173 = U284/U237/vout (480 , -694)
*       173 = U284/U238/B (494.5 , -677.5)
*       175 = U284/Carry (602.5 , -707.5)
*       175 = U249/U210/A (549 , -745.5)
*       175 = U249/AA (549 , -739.5)
*       175 = U284/U238/C (602.5 , -675)
*       177 = U249/U210/B (455.5 , -747.5)
*       177 = U249/BB (455.5 , -739)
*       177 = U249/U229/vout (414 , -761)
*       181 = U247/U210/C (279.5 , -745)
*       181 = U247/U213/A (316 , -747)
*       182 = U247/U210/A (265 , -745.5)
*       182 = U247/AA (265 , -739.5)
*       182 = U283/Carry (318.5 , -707.5)
*       182 = U283/U238/C (318.5 , -675)
*       187 = U247/U210/B (171.5 , -747.5)
*       187 = U247/BB (171.5 , -739)
*       187 = U247/U229/vout (130 , -761)
*       188 = U283/Sum (202.5 , -708)
*       188 = U249/CC (474.5 , -739)
*       188 = U249/U211/A (549 , -796.5)
*       188 = U283/U238/S (202.5 , -677)
*       189 = U283/U237/vout (196 , -694)
*       189 = U283/U238/B (210.5 , -677.5)
*       192 = U282/Sum (-82 , -708)
*       192 = U247/CC (190.5 , -739)
*       192 = U247/U211/A (265 , -796.5)
*       192 = U282/U238/S (-82 , -677)
*       196 = U245/U210/C (-5 , -745)
*       196 = U245/U213/A (31.5 , -747)
*       197 = U245/U210/A (-19.5 , -745.5)
*       197 = U245/AA (-19.5 , -739.5)
*       197 = U282/Carry (34 , -707.5)
*       197 = U282/U238/C (34 , -675)
*       201 = U245/U210/B (-113 , -747.5)
*       201 = U245/BB (-113 , -739)
*       201 = U245/U229/vout (-154.5 , -761)
*       202 = U282/U238/B (-74 , -677.5)
*       202 = U282/U237/vout (-88.5 , -694)
*       203 = U279/U215/vin (-235.5 , -717.5)
*       203 = U279/U213/O/P (-224 , -659)
*       214 = U243/U210/A (-304 , -745.5)
*       214 = U243/AA (-304 , -739.5)
*       214 = U279/U215/vout (-250 , -716)
*       214 = U279/Carry (-250.5 , -731)
*       215 = U279/U211/C (-289.5 , -700)
*       215 = U279/U213/B (-237.5 , -652.5)
*       216 = U243/U210/C (-289.5 , -745)
*       216 = U243/U213/A (-253 , -747)
*       219 = U243/U210/B (-397.5 , -747.5)
*       219 = U243/BB (-397.5 , -739)
*       219 = U243/U229/vout (-439 , -761)
*       220 = U279/Sum (-405.5 , -731.5)
*       220 = U245/CC (-94 , -739)
*       220 = U245/U211/A (-19.5 , -796.5)
*       220 = U279/U211/S (-405.5 , -702)
*       221 = U279/U228/OUTPUT (-425 , -709.5)
*       221 = U279/U229/vin (-424.5 , -666.5)
*       222 = U279/U211/B (-397.5 , -702.5)
*       222 = U279/U210/S (-405.5 , -651)
*       224 = U241/U213/A (-537.5 , -747)
*       224 = U241/U210/C (-574 , -745)
*       228 = U281/U238/S (-663.5 , -678)
*       228 = U281/Sum (-663.5 , -709)
*       228 = U243/U211/A (-304 , -796.5)
*       228 = U243/CC (-378.5 , -739)
*       232 = U241/U210/A (-588.5 , -745.5)
*       232 = U241/AA (-588.5 , -739.5)
*       232 = U281/Carry (-547.5 , -708.5)
*       232 = U281/U238/C (-547.5 , -676)
*       234 = U241/U229/vout (-723.5 , -761)
*       234 = U241/U210/B (-682 , -747.5)
*       234 = U241/BB (-682 , -739)
*       235 = U281/U237/vin (-698.5 , -694)
*       235 = U281/U234/OUTPUT (-709.5 , -685.5)
*       236 = U241/U210/S (-690 , -747)
*       236 = U241/U211/B (-682 , -798.5)
*       238 = U299/U232/S (-976.4 , -677.9)
*       238 = U299/Sum (-976.5 , -708)
*       238 = U241/CC (-663 , -739)
*       238 = U241/U211/A (-588.5 , -796.5)
*       242 = U299/U232/A (-874.9 , -676.4)
*       242 = U299/AA (-875 , -671.5)
*       242 = U298/Carry (-860 , -629.5)
*       242 = U298/U232/C (-860.4 , -597.9)
*       244 = U300/U232/A (-874.9 , -771.4)
*       244 = U300/AA (-875 , -766.5)
*       244 = U299/Carry (-860 , -707.5)
*       244 = U299/U232/C (-860.4 , -675.9)
*       245 = U300/U232/B (-968.4 , -773.4)
*       245 = U300/U234/OUTPUT (-986.5 , -780.5)
*       247 = U326/DataInB (-1557.5 , -715)
*       248 = U326/DataIn (-1557.5 , -739)
*       248 = U300/U234/INPUTA (-1067 , -798)
*       248 = U300/X (-1072 , -784)
*       248 = X2 (-1073 , -786.5)
*       248 = U241/X (-795 , -784)
*       248 = U241/U228/INPUTA (-790 , -823)
*       248 = U243/U228/INPUTA (-505.5 , -823)
*       248 = U243/X (-510.5 , -784)
*       248 = U245/U228/INPUTA (-221 , -823)
*       248 = U245/X (-226 , -784)
*       248 = U247/U228/INPUTA (63.5 , -823)
*       248 = U247/X (58.5 , -784)
*       248 = U249/U228/INPUTA (347.5 , -823)
*       248 = U249/X (342.5 , -784)
*       248 = U251/U228/INPUTA (632 , -823)
*       248 = U251/X (627 , -784)
*       249 = U326/DataInUnBuf (-1557.5 , -699)
*       250 = U252/U213/A (884.5 , -843)
*       250 = U252/U210/C (848 , -841)
*       251 = U251/U215/vin (902 , -813.5)
*       251 = U251/U213/O/P (913.5 , -755)
*       252 = U251/U213/B (900 , -748.5)
*       252 = U251/U211/C (848 , -796)
*       263 = U251/U211/B (740 , -798.5)
*       263 = U251/U210/S (732 , -747)
*       265 = U251/Sum (732 , -827.5)
*       265 = U251/U211/S (732 , -798)
*       265 = P2 (922 , -800.5)
*       265 = U341/DataOut (1494.5 , -1041)
*       267 = U252/U210/A (833.5 , -841.5)
*       267 = U252/AA (833.5 , -835.5)
*       267 = U251/U215/vout (887.5 , -812)
*       267 = U251/Carry (887 , -827)
*       268 = U252/U229/vout (698.5 , -857)
*       268 = U252/U210/B (740 , -843.5)
*       268 = U252/BB (740 , -835)
*       269 = U252/U229/vin (713 , -858.5)
*       269 = U252/U228/OUTPUT (712.5 , -901.5)
*       272 = U249/U215/vin (617.5 , -813.5)
*       272 = U249/U213/O/P (629 , -755)
*       273 = U250/U213/A (600 , -843)
*       273 = U250/U210/C (563.5 , -841)
*       274 = U249/U211/C (563.5 , -796)
*       274 = U249/U213/B (615.5 , -748.5)
*       283 = U249/U211/B (455.5 , -798.5)
*       283 = U249/U210/S (447.5 , -747)
*       285 = U249/Sum (447.5 , -827.5)
*       285 = U252/CC (759 , -835)
*       285 = U252/U211/A (833.5 , -892.5)
*       285 = U249/U211/S (447.5 , -798)
*       288 = U250/U210/A (549 , -841.5)
*       288 = U250/AA (549 , -835.5)
*       288 = U249/U215/vout (603 , -812)
*       288 = U249/Carry (602.5 , -827)
*       290 = U249/U228/OUTPUT (428 , -805.5)
*       290 = U249/U229/vin (428.5 , -762.5)
*       291 = U247/U215/vin (333.5 , -813.5)
*       291 = U247/U213/O/P (345 , -755)
*       292 = U250/U210/B (455.5 , -843.5)
*       292 = U250/BB (455.5 , -835)
*       292 = U250/U229/vout (414 , -857)
*       295 = U248/U210/A (265 , -841.5)
*       295 = U248/AA (265 , -835.5)
*       295 = U247/U215/vout (319 , -812)
*       295 = U247/Carry (318.5 , -827)
*       296 = U248/U210/C (279.5 , -841)
*       296 = U248/U213/A (316 , -843)
*       297 = U247/U211/C (279.5 , -796)
*       297 = U247/U213/B (331.5 , -748.5)
*       305 = U248/U210/B (171.5 , -843.5)
*       305 = U248/BB (171.5 , -835)
*       305 = U248/U229/vout (130 , -857)
*       307 = U247/U228/OUTPUT (144 , -805.5)
*       307 = U247/U229/vin (144.5 , -762.5)
*       308 = U247/U211/B (171.5 , -798.5)
*       308 = U247/U210/S (163.5 , -747)
*       310 = U247/Sum (163.5 , -827.5)
*       310 = U247/U211/S (163.5 , -798)
*       310 = U250/CC (474.5 , -835)
*       310 = U250/U211/A (549 , -892.5)
*       313 = U245/U215/vin (49 , -813.5)
*       313 = U245/U213/O/P (60.5 , -755)
*       320 = U246/U210/A (-19.5 , -841.5)
*       320 = U246/AA (-19.5 , -835.5)
*       320 = U245/U215/vout (34.5 , -812)
*       320 = U245/Carry (34 , -827)
*       321 = U246/U210/C (-5 , -841)
*       321 = U246/U213/A (31.5 , -843)
*       322 = U245/U211/C (-5 , -796)
*       322 = U245/U213/B (47 , -748.5)
*       328 = U246/U210/B (-113 , -843.5)
*       328 = U246/BB (-113 , -835)
*       328 = U246/U229/vout (-154.5 , -857)
*       329 = U245/Sum (-121 , -827.5)
*       329 = U248/CC (190.5 , -835)
*       329 = U248/U211/A (265 , -892.5)
*       329 = U245/U211/S (-121 , -798)
*       330 = U245/U228/OUTPUT (-140.5 , -805.5)
*       330 = U245/U229/vin (-140 , -762.5)
*       331 = U245/U211/B (-113 , -798.5)
*       331 = U245/U210/S (-121 , -747)
*       334 = U308/U228/INPUTB (-165.5 , -962)
*       334 = U246/U228/INPUTB (-165.5 , -917)
*       334 = U246/Y (-164 , -836.5)
*       334 = U245/U228/INPUTB (-165.5 , -821)
*       334 = U245/Y (-164 , -740.5)
*       334 = U288/U239/B (-150.5 , -615)
*       334 = U282/U234/INPUTB (-153 , -700)
*       334 = U282/Y (-151 , -671)
*       334 = U288/Y (-151 , -591)
*       334 = Y3 (-151 , -591)
*       334 = U317/DataIn (-126.5 , 446)
*       335 = U243/U215/vin (-235.5 , -813.5)
*       335 = U243/U213/O/P (-224 , -755)
*       344 = U244/U210/A (-304 , -841.5)
*       344 = U244/AA (-304 , -835.5)
*       344 = U243/U215/vout (-250 , -812)
*       344 = U243/Carry (-250.5 , -827)
*       345 = U244/U210/C (-289.5 , -841)
*       345 = U244/U213/A (-253 , -843)
*       346 = U243/U211/C (-289.5 , -796)
*       346 = U243/U213/B (-237.5 , -748.5)
*       351 = U244/U210/B (-397.5 , -843.5)
*       351 = U244/BB (-397.5 , -835)
*       351 = U244/U229/vout (-439 , -857)
*       352 = U243/U228/OUTPUT (-425 , -805.5)
*       352 = U243/U229/vin (-424.5 , -762.5)
*       353 = U243/U211/B (-397.5 , -798.5)
*       353 = U243/U210/S (-405.5 , -747)
*       354 = U243/Sum (-405.5 , -827.5)
*       354 = U243/U211/S (-405.5 , -798)
*       354 = U246/CC (-94 , -835)
*       354 = U246/U211/A (-19.5 , -892.5)
*       356 = U242/U213/A (-537.5 , -843)
*       356 = U242/U210/C (-574 , -841)
*       357 = U241/U215/vin (-520 , -813.5)
*       357 = U241/U213/O/P (-508.5 , -755)
*       358 = U241/U213/B (-522 , -748.5)
*       358 = U241/U211/C (-574 , -796)
*       367 = U242/U210/A (-588.5 , -841.5)
*       367 = U242/AA (-588.5 , -835.5)
*       367 = U241/U215/vout (-534.5 , -812)
*       367 = U241/Carry (-535 , -827)
*       372 = U242/U229/vout (-723.5 , -857)
*       372 = U242/U210/B (-682 , -843.5)
*       372 = U242/BB (-682 , -835)
*       373 = U241/Sum (-690 , -827.5)
*       373 = U244/U211/A (-304 , -892.5)
*       373 = U244/CC (-378.5 , -835)
*       373 = U241/U211/S (-690 , -798)
*       374 = U242/U210/S (-690 , -843)
*       374 = U242/U211/B (-682 , -894.5)
*       375 = U241/U228/OUTPUT (-709.5 , -805.5)
*       375 = U241/U229/vin (-709 , -762.5)
*       381 = U242/CC (-663 , -835)
*       381 = U242/U211/A (-588.5 , -892.5)
*       381 = U300/U232/S (-976.4 , -772.9)
*       381 = U300/Sum (-976.5 , -803)
*       383 = U301/U232/A (-874.9 , -867.4)
*       383 = U301/AA (-875 , -862.5)
*       383 = U300/U232/C (-860.4 , -770.9)
*       383 = U300/Carry (-860 , -802.5)
*       384 = U301/U232/B (-968.4 , -869.4)
*       384 = U301/U234/OUTPUT (-986.5 , -876.5)
*       388 = U294/U213/A (875 , -939)
*       388 = U294/U210/C (838.5 , -937)
*       389 = U252/U215/vin (902 , -909.5)
*       389 = U252/U213/O/P (913.5 , -851)
*       390 = U252/U213/B (900 , -844.5)
*       390 = U252/U211/C (848 , -892)
*       402 = U252/U211/B (740 , -894.5)
*       402 = U252/U210/S (732 , -843)
*       403 = U252/Sum (732 , -923.5)
*       403 = U252/U211/S (732 , -894)
*       403 = P3 (922 , -896.5)
*       403 = U340/DataOut (1494.5 , -1477)
*       404 = U294/U210/A (824 , -937.5)
*       404 = U294/AA (824 , -931.5)
*       404 = U252/U215/vout (887.5 , -908)
*       404 = U252/Carry (887 , -923)
*       405 = U294/U210/B (730.5 , -939.5)
*       405 = U294/BB (730.5 , -931)
*       405 = U294/U228/OUTPUT (712.5 , -946.5)
*       408 = U250/U215/vin (617.5 , -909.5)
*       408 = U250/U213/O/P (629 , -851)
*       409 = U295/U213/A (590.5 , -939)
*       409 = U295/U210/C (554 , -937)
*       410 = U250/U211/C (563.5 , -892)
*       410 = U250/U213/B (615.5 , -844.5)
*       420 = U250/Sum (447.5 , -923.5)
*       420 = U294/CC (749.5 , -931)
*       420 = U294/U211/A (824 , -988.5)
*       420 = U250/U211/S (447.5 , -894)
*       423 = U250/U211/B (455.5 , -894.5)
*       423 = U250/U210/S (447.5 , -843)
*       425 = U295/U210/A (539.5 , -937.5)
*       425 = U295/AA (539.5 , -931.5)
*       425 = U250/U215/vout (603 , -908)
*       425 = U250/Carry (602.5 , -923)
*       427 = U248/Sum (163.5 , -923.5)
*       427 = U295/CC (465 , -931)
*       427 = U295/U211/A (539.5 , -988.5)
*       427 = U248/U211/S (163.5 , -894)
*       428 = U295/U210/B (446 , -939.5)
*       428 = U295/BB (446 , -931)
*       428 = U295/U228/OUTPUT (428 , -946.5)
*       429 = U250/U229/vin (428.5 , -858.5)
*       429 = U250/U228/OUTPUT (428 , -901.5)
*       430 = U248/U215/vin (333.5 , -909.5)
*       430 = U248/U213/O/P (345 , -851)
*       433 = U297/U213/A (306.5 , -939)
*       433 = U297/U210/C (270 , -937)
*       434 = U248/U211/C (279.5 , -892)
*       434 = U248/U213/B (331.5 , -844.5)
*       439 = U248/U229/vin (144.5 , -858.5)
*       439 = U248/U228/OUTPUT (144 , -901.5)
*       441 = U248/U211/B (171.5 , -894.5)
*       441 = U248/U210/S (163.5 , -843)
*       442 = U325/DataIn (-1557.5 , -1175)
*       442 = U301/U234/INPUTA (-1067 , -894)
*       442 = U301/X (-1072 , -880)
*       442 = X3 (-1073 , -882.5)
*       442 = U242/X (-795 , -880)
*       442 = U242/U228/INPUTA (-790 , -919)
*       442 = U244/U228/INPUTA (-505.5 , -919)
*       442 = U244/X (-510.5 , -880)
*       442 = U246/U228/INPUTA (-221 , -919)
*       442 = U246/X (-226 , -880)
*       442 = U248/U228/INPUTA (63.5 , -919)
*       442 = U248/X (58.5 , -880)
*       442 = U250/U228/INPUTA (347.5 , -919)
*       442 = U250/X (342.5 , -880)
*       442 = U252/U228/INPUTA (632 , -919)
*       442 = U252/X (627 , -880)
*       445 = U297/U210/A (255.5 , -937.5)
*       445 = U297/AA (255.5 , -931.5)
*       445 = U248/U215/vout (319 , -908)
*       445 = U248/Carry (318.5 , -923)
*       451 = U297/U210/B (162 , -939.5)
*       451 = U297/BB (162 , -931)
*       451 = U297/U228/OUTPUT (144 , -946.5)
*       452 = U246/U215/vin (49 , -909.5)
*       452 = U246/U213/O/P (60.5 , -851)
*       457 = U308/U210/A (-29 , -937.5)
*       457 = U308/AA (-29 , -931.5)
*       457 = U246/U215/vout (34.5 , -908)
*       457 = U246/Carry (34 , -923)
*       458 = U308/U210/C (-14.5 , -937)
*       458 = U308/U213/A (22 , -939)
*       459 = U246/U211/C (-5 , -892)
*       459 = U246/U213/B (47 , -844.5)
*       467 = U246/Sum (-121 , -923.5)
*       467 = U297/CC (181 , -931)
*       467 = U297/U211/A (255.5 , -988.5)
*       467 = U246/U211/S (-121 , -894)
*       468 = U246/U229/vin (-140 , -858.5)
*       468 = U246/U228/OUTPUT (-140.5 , -901.5)
*       469 = U246/U211/B (-113 , -894.5)
*       469 = U246/U210/S (-121 , -843)
*       472 = U308/U210/B (-122.5 , -939.5)
*       472 = U308/BB (-122.5 , -931)
*       472 = U308/U228/OUTPUT (-140.5 , -946.5)
*       473 = U244/U215/vin (-235.5 , -909.5)
*       473 = U244/U213/O/P (-224 , -851)
*       481 = U309/U210/A (-313.5 , -937.5)
*       481 = U309/AA (-313.5 , -931.5)
*       481 = U244/U215/vout (-250 , -908)
*       481 = U244/Carry (-250.5 , -923)
*       482 = U309/U210/C (-299 , -937)
*       482 = U309/U213/A (-262.5 , -939)
*       483 = U244/U211/C (-289.5 , -892)
*       483 = U244/U213/B (-237.5 , -844.5)
*       488 = U244/U229/vin (-424.5 , -858.5)
*       488 = U244/U228/OUTPUT (-425 , -901.5)
*       489 = U244/U211/B (-397.5 , -894.5)
*       489 = U244/U210/S (-405.5 , -843)
*       490 = U244/Sum (-405.5 , -923.5)
*       490 = U244/U211/S (-405.5 , -894)
*       490 = U308/CC (-103.5 , -931)
*       490 = U308/U211/A (-29 , -988.5)
*       493 = U309/U210/B (-407 , -939.5)
*       493 = U309/BB (-407 , -931)
*       493 = U309/U228/OUTPUT (-425 , -946.5)
*       494 = U242/U215/vin (-520 , -909.5)
*       494 = U242/U213/O/P (-508.5 , -851)
*       495 = U242/U213/B (-522 , -844.5)
*       495 = U242/U211/C (-574 , -892)
*       499 = U310/U213/B (-531.5 , -940.5)
*       499 = U310/U211/C (-583.5 , -988)
*       502 = U310/U213/A (-547 , -939)
*       502 = U310/U210/C (-583.5 , -937)
*       507 = U310/U210/A (-598 , -937.5)
*       507 = U310/AA (-598 , -931.5)
*       507 = U242/U215/vout (-534.5 , -908)
*       507 = U242/Carry (-535 , -923)
*       510 = U310/U210/B (-691.5 , -939.5)
*       510 = U310/BB (-691.5 , -931)
*       510 = U310/U228/OUTPUT (-709.5 , -946.5)
*       511 = U242/Sum (-690 , -923.5)
*       511 = U309/U211/A (-313.5 , -988.5)
*       511 = U309/CC (-388 , -931)
*       511 = U242/U211/S (-690 , -894)
*       512 = U242/U229/vin (-709 , -858.5)
*       512 = U242/U228/OUTPUT (-709.5 , -901.5)
*       516 = U302/U238/A (-839 , -962.5)
*       516 = U302/AA (-839 , -958.5)
*       516 = U301/U232/C (-860.4 , -866.9)
*       516 = U301/Carry (-860 , -898.5)
*       520 = U302/U237/vout (-947 , -981)
*       520 = U302/U238/B (-932.5 , -964.5)
*       521 = U302/U238/S (-940.5 , -964)
*       521 = U302/Sum (-940.5 , -995)
*       521 = U304/U210/B (-691.5 , -1041.5)
*       521 = U304/BB (-691.5 , -1033)
*       522 = U310/U211/A (-598 , -988.5)
*       522 = U310/CC (-672.5 , -931)
*       522 = U301/U232/S (-976.4 , -868.9)
*       522 = U301/Sum (-976.5 , -899)
*       524 = U302/U237/vin (-975.5 , -980)
*       524 = U302/U234/OUTPUT (-986.5 , -971.5)
*       528 = U294/U213/B (890.5 , -940.5)
*       528 = U294/U211/C (838.5 , -988)
*       530 = U294/U215/vin (892.5 , -1005.5)
*       530 = U294/U213/O/P (904 , -947)
*       536 = U269/S (722.5 , -1041)
*       536 = P5 (912.5 , -1045.5)
*       536 = U337/DataOut (1319.5 , -2174)
*       537 = U294/Sum (722.5 , -1019.5)
*       537 = U294/U211/S (722.5 , -990)
*       537 = P4 (912.5 , -992.5)
*       537 = U339/DataOut (1494.5 , -1913)
*       539 = U294/U211/B (730.5 , -990.5)
*       539 = U294/U210/S (722.5 , -939)
*       541 = U294/Carry (877.5 , -1019)
*       541 = U269/A (824 , -1039.5)
*       541 = U294/U215/vout (878 , -1004)
*       542 = U296/U213/A (590.5 , -1041)
*       542 = U296/U210/C (554 , -1039)
*       543 = U295/U213/B (606 , -940.5)
*       543 = U295/U211/C (554 , -988)
*       545 = U295/U215/vin (608 , -1005.5)
*       545 = U295/U213/O/P (619.5 , -947)
*       554 = U295/Sum (438 , -1019.5)
*       554 = U269/B (730.5 , -1041.5)
*       554 = U295/U211/S (438 , -990)
*       556 = U295/U211/B (446 , -990.5)
*       556 = U295/U210/S (438 , -939)
*       558 = U296/U210/A (539.5 , -1039.5)
*       558 = U296/AA (539.5 , -1033.5)
*       558 = U295/Carry (593 , -1019)
*       558 = U295/U215/vout (593.5 , -1004)
*       559 = U296/CC (465 , -1033)
*       559 = U296/U211/A (539.5 , -1090.5)
*       559 = U269/C (838.5 , -1039)
*       560 = U297/U215/vin (324 , -1005.5)
*       560 = U297/U213/O/P (335.5 , -947)
*       562 = U307/U213/A (306.5 , -1041)
*       562 = U307/U210/C (270 , -1039)
*       563 = U297/U211/C (270 , -988)
*       563 = U297/U213/B (322 , -940.5)
*       566 = U297/Sum (154 , -1019.5)
*       566 = U296/U210/B (446 , -1041.5)
*       566 = U296/BB (446 , -1033)
*       566 = U297/U211/S (154 , -990)
*       568 = U307/CC (181 , -1033)
*       568 = U307/U211/A (255.5 , -1090.5)
*       568 = U296/U215/vout (593.5 , -1106)
*       568 = U296/Carry (593 , -1121)
*       569 = U297/U211/B (162 , -990.5)
*       569 = U297/U210/S (154 , -939)
*       573 = U307/U210/A (255.5 , -1039.5)
*       573 = U307/AA (255.5 , -1033.5)
*       573 = U297/Carry (309 , -1019)
*       573 = U297/U215/vout (309.5 , -1004)
*       577 = U308/U215/vin (39.5 , -1005.5)
*       577 = U308/U213/O/P (51 , -947)
*       580 = U306/U210/A (-29 , -1039.5)
*       580 = U306/AA (-29 , -1033.5)
*       580 = U308/Carry (24.5 , -1019)
*       580 = U308/U215/vout (25 , -1004)
*       581 = U308/U211/C (-14.5 , -988)
*       581 = U308/U213/B (37.5 , -940.5)
*       583 = U306/U210/C (-14.5 , -1039)
*       583 = U306/U213/A (22 , -1041)
*       592 = U308/Sum (-130.5 , -1019.5)
*       592 = U307/U210/B (162 , -1041.5)
*       592 = U307/BB (162 , -1033)
*       592 = U308/U211/S (-130.5 , -990)
*       593 = U306/CC (-103.5 , -1033)
*       593 = U306/U211/A (-29 , -1090.5)
*       593 = U307/U215/vout (309.5 , -1106)
*       593 = U307/Carry (309 , -1121)
*       594 = U308/U211/B (-122.5 , -990.5)
*       594 = U308/U210/S (-130.5 , -939)
*       595 = U309/U215/vin (-245 , -1005.5)
*       595 = U309/U213/O/P (-233.5 , -947)
*       602 = U305/U210/A (-313.5 , -1039.5)
*       602 = U305/AA (-313.5 , -1033.5)
*       602 = U309/Carry (-260 , -1019)
*       602 = U309/U215/vout (-259.5 , -1004)
*       603 = U309/U211/C (-299 , -988)
*       603 = U309/U213/B (-247 , -940.5)
*       604 = U305/U210/C (-299 , -1039)
*       604 = U305/U213/A (-262.5 , -1041)
*       610 = U309/Sum (-415 , -1019.5)
*       610 = U306/U210/B (-122.5 , -1041.5)
*       610 = U306/BB (-122.5 , -1033)
*       610 = U309/U211/S (-415 , -990)
*       611 = U305/U211/A (-313.5 , -1090.5)
*       611 = U305/CC (-388 , -1033)
*       611 = U306/U215/vout (25 , -1106)
*       611 = U306/Carry (24.5 , -1121)
*       612 = U309/U211/B (-407 , -990.5)
*       612 = U309/U210/S (-415 , -939)
*       613 = U310/U215/vin (-529.5 , -1005.5)
*       613 = U310/U213/O/P (-518 , -947)
*       618 = U304/U213/B (-531.5 , -1042.5)
*       618 = U304/U211/C (-583.5 , -1090)
*       621 = U304/U213/A (-547 , -1041)
*       621 = U304/U210/C (-583.5 , -1039)
*       624 = U304/U210/A (-598 , -1039.5)
*       624 = U304/AA (-598 , -1033.5)
*       624 = U310/Carry (-544.5 , -1019)
*       624 = U310/U215/vout (-544 , -1004)
*       628 = U310/Sum (-699.5 , -1019.5)
*       628 = U305/U210/B (-407 , -1041.5)
*       628 = U305/BB (-407 , -1033)
*       628 = U310/U211/S (-699.5 , -990)
*       629 = U310/U211/B (-691.5 , -990.5)
*       629 = U310/U210/S (-699.5 , -939)
*       630 = U303/U213/A (-844.5 , -1041)
*       630 = U303/U210/C (-881 , -1039)
*       639 = U303/U210/A (-895.5 , -1039.5)
*       639 = U303/AA (-895.5 , -1033.5)
*       639 = U304/U215/vout (-544 , -1106)
*       639 = U304/Carry (-544.5 , -1121)
*       645 = U296/U215/vin (608 , -1107.5)
*       645 = U296/U213/O/P (619.5 , -1049)
*       646 = U296/U213/B (606 , -1042.5)
*       646 = U296/U211/C (554 , -1090)
*       650 = U296/U211/B (446 , -1092.5)
*       650 = U296/U210/S (438 , -1041)
*       651 = U307/U215/vin (324 , -1107.5)
*       651 = U307/U213/O/P (335.5 , -1049)
*       652 = U307/U211/C (270 , -1090)
*       652 = U307/U213/B (322 , -1042.5)
*       655 = U307/U211/B (162 , -1092.5)
*       655 = U307/U210/S (154 , -1041)
*       657 = U306/U215/vin (39.5 , -1107.5)
*       657 = U306/U213/O/P (51 , -1049)
*       659 = U306/U211/C (-14.5 , -1090)
*       659 = U306/U213/B (37.5 , -1042.5)
*       662 = U306/U211/B (-122.5 , -1092.5)
*       662 = U306/U210/S (-130.5 , -1041)
*       663 = U305/U215/vin (-245 , -1107.5)
*       663 = U305/U213/O/P (-233.5 , -1049)
*       666 = U305/U211/C (-299 , -1090)
*       666 = U305/U213/B (-247 , -1042.5)
*       668 = U305/U211/B (-407 , -1092.5)
*       668 = U305/U210/S (-415 , -1041)
*       669 = U304/U215/vin (-529.5 , -1107.5)
*       669 = U304/U213/O/P (-518 , -1049)
*       673 = U304/U211/A (-598 , -1090.5)
*       673 = U304/CC (-672.5 , -1033)
*       673 = U305/U215/vout (-259.5 , -1106)
*       673 = U305/Carry (-260 , -1121)
*       674 = U304/U211/B (-691.5 , -1092.5)
*       674 = U304/U210/S (-699.5 , -1041)
*       675 = U303/U215/vin (-827 , -1107.5)
*       675 = U303/U213/O/P (-815.5 , -1049)
*       676 = U303/U215/vout (-841.5 , -1106)
*       676 = U303/Carry (-842 , -1121)
*       677 = U303/U213/B (-829 , -1042.5)
*       677 = U303/U211/C (-881 , -1090)
*       681 = U303/U211/B (-989 , -1092.5)
*       681 = U303/U210/S (-997 , -1041)
*       682 = U303/U211/A (-895.5 , -1090.5)
*       682 = U303/CC (-970 , -1033)
*       682 = U302/U238/C (-824.5 , -962)
*       682 = U302/Carry (-824.5 , -994.5)
*       683 = U325/DataInB (-1557.5 , -1151)
*       684 = U325/DataInUnBuf (-1557.5 , -1135)
*       687 = U334/DataOut (11.5 , -2174)
*       687 = U306/Sum (-130.5 , -1121.5)
*       687 = P8 (-130.5 , -1123)
*       687 = U306/U211/S (-130.5 , -1092)
*       688 = U324/DataInUnBuf (-1557.5 , -1571)
*       696 = U324/DataIn (-1557.5 , -1611)
*       696 = U302/U234/INPUTA (-1067 , -989)
*       696 = U302/X (-1072 , -975.5)
*       696 = X4 (-1073 , -977.5)
*       696 = U310/U228/INPUTA (-790 , -964)
*       696 = U310/X (-795 , -976)
*       696 = U309/U228/INPUTA (-505.5 , -964)
*       696 = U309/X (-510.5 , -976)
*       696 = U308/U228/INPUTA (-221 , -964)
*       696 = U308/X (-226 , -976)
*       696 = U297/U228/INPUTA (63.5 , -964)
*       696 = U297/X (58.5 , -976)
*       696 = U295/U228/INPUTA (347.5 , -964)
*       696 = U295/X (342.5 , -976)
*       696 = U294/U228/INPUTA (632 , -964)
*       696 = U294/X (627 , -976)
*       697 = U324/DataInB (-1557.5 , -1587)
*       698 = U336/DataOut (883.5 , -2174)
*       698 = U296/Sum (438 , -1121.5)
*       698 = P6 (438 , -1123)
*       698 = U296/U211/S (438 , -1092)
*       699 = U335/DataOut (447.5 , -2174)
*       699 = U307/Sum (154 , -1121.5)
*       699 = P7 (154 , -1123)
*       699 = U307/U211/S (154 , -1092)
*       734 = U333/DataOut (-424.5 , -2174)
*       734 = U305/Sum (-415 , -1121.5)
*       734 = P9 (-415 , -1123)
*       734 = U305/U211/S (-415 , -1092)
*       741 = U332/DataOut (-860.5 , -2174)
*       741 = U304/Sum (-699.5 , -1121.5)
*       741 = P10 (-699.5 , -1123)
*       741 = U304/U211/S (-699.5 , -1092)
*       747 = U330/DataOut (-1296.5 , -2174)
*       747 = U303/Sum (-997 , -1121.5)
*       747 = P11 (-997 , -1123)
*       747 = U303/U211/S (-997 , -1092)


Cpar1 1 0 643.3195f
Cpar2 2 0 643.3195f
Cpar3 3 0 643.3195f
Cpar4 4 0 643.3195f
Cpar5 5 0 643.3195f
Cpar6 6 0 643.3195f
Cpar7 7 0 643.3195f
Cpar8 8 0 48.635973p
Cpar9 9 0 20.365125f
Cpar10 10 0 74.2155f
Cpar11 11 0 44.412313f
Cpar12 12 0 76.08327p
Cpar13 13 0 44.412313f
Cpar14 14 0 20.365125f
Cpar15 15 0 44.412313f
Cpar16 16 0 20.365125f
Cpar17 17 0 30.276625f
Cpar18 18 0 126.67555f
Cpar19 19 0 20.365125f
Cpar20 20 0 74.2155f
Cpar21 21 0 44.412313f
Cpar22 22 0 44.412313f
Cpar23 23 0 20.365125f
Cpar24 24 0 30.276625f
Cpar25 25 0 44.412313f
Cpar26 26 0 20.365125f
Cpar27 27 0 74.2155f
Cpar28 28 0 20.365125f
Cpar29 29 0 74.2155f
Cpar30 30 0 44.412313f
Cpar31 31 0 30.276625f
Cpar32 32 0 74.2155f
Cpar33 33 0 30.276625f
Cpar34 34 0 74.2155f
Cpar35 35 0 30.276625f
Cpar36 36 0 74.2155f
Cpar37 37 0 126.72528f
Cpar38 38 0 30.276625f
Cpar39 39 0 30.276625f
Cpar40 40 0 126.73794f
Cpar41 41 0 127.54375f
Cpar42 42 0 74.2155f
Cpar43 43 0 44.412313f
Cpar44 44 0 20.365125f
Cpar45 45 0 130.79081f
Cpar46 46 0 30.276625f
Cpar47 47 0 643.3195f
Cpar48 48 0 643.3195f
Cpar49 49 0 74.2155f
Cpar50 50 0 74.2155f
Cpar51 51 0 30.276625f
Cpar52 52 0 44.412313f
Cpar53 53 0 20.365125f
Cpar54 54 0 132.30608f
Cpar55 55 0 20.365125f
Cpar56 56 0 44.412312f
Cpar57 57 0 120.49825f
Cpar58 58 0 30.276625f
Cpar59 59 0 643.3195f
Cpar60 60 0 643.3195f
Cpar61 61 0 74.2155f
Cpar62 62 0 3.8650312f
Cpar63 63 0 44.412313f
Cpar64 64 0 20.365125f
Cpar65 65 0 3.7905312f
Cpar66 67 0 2.52975f
Cpar67 68 0 4.0961875f
Cpar68 69 0 3.24375f
Cpar69 70 0 3.3804063f
Cpar70 71 0 12.825703f
Cpar71 72 0 8.3536875f
Cpar72 73 0 127.11641f
Cpar73 76 0 3.7905312f
Cpar74 77 0 2.52975f
Cpar75 78 0 4.0961875f
Cpar76 80 0 3.24375f
Cpar77 82 0 4.8002188f
Cpar78 83 0 126.80463f
Cpar79 84 0 3.3804063f
Cpar80 85 0 12.825703f
Cpar81 88 0 3.7905312f
Cpar82 89 0 2.52975f
Cpar83 90 0 4.0961875f
Cpar84 91 0 3.3804063f
Cpar85 94 0 4.8139688f
Cpar86 95 0 12.825703f
Cpar87 97 0 2.52975f
Cpar88 98 0 4.0961875f
Cpar89 99 0 3.7905312f
Cpar90 100 0 3.24375f
Cpar91 101 0 3.3804063f
Cpar92 104 0 4.8002188f
Cpar93 105 0 12.825703f
Cpar94 107 0 1.04175f
Cpar95 108 0 3.2747812f
Cpar96 110 0 2.52975f
Cpar97 111 0 3.7905312f
Cpar98 112 0 2.52975f
Cpar99 113 0 4.0961875f
Cpar100 114 0 3.2903437f
Cpar101 115 0 4.0961875f
Cpar102 116 0 23.349219f
Cpar103 117 0 3.24375f
Cpar104 118 0 3.7905312f
Cpar105 119 0 3.24375f
Cpar106 120 0 3.6394063f
Cpar107 121 0 12.825703f
Cpar108 124 0 2.52975f
Cpar109 125 0 4.0961875f
Cpar110 126 0 3.7905312f
Cpar111 127 0 3.24375f
Cpar112 128 0 3.3804063f
Cpar113 130 0 3.8650313f
Cpar114 132 0 4.7388906f
Cpar115 135 0 2.52975f
Cpar116 136 0 4.0961875f
Cpar117 137 0 3.7905312f
Cpar118 138 0 2.52975f
Cpar119 139 0 4.0961875f
Cpar120 140 0 3.7905312f
Cpar121 141 0 3.24375f
Cpar122 142 0 3.24375f
Cpar123 143 0 23.378487f
Cpar124 144 0 12.806188f
Cpar125 146 0 12.806188f
Cpar126 148 0 44.412313f
Cpar127 149 0 20.365125f
Cpar128 150 0 74.2155f
Cpar129 151 0 30.276625f
Cpar130 152 0 120.49825f
Cpar131 153 0 3.2903437f
Cpar132 156 0 1.04175f
Cpar133 157 0 2.52975f
Cpar134 158 0 4.0961875f
Cpar135 159 0 3.7905312f
Cpar136 160 0 25.727406f
Cpar137 161 0 3.8650312f
Cpar138 162 0 3.24375f
Cpar139 163 0 3.3376875f
Cpar140 164 0 3.6394063f
Cpar141 165 0 12.786219f
Cpar142 166 0 1.04175f
Cpar143 167 0 3.2903437f
Cpar144 170 0 2.52975f
Cpar145 171 0 4.0961875f
Cpar146 172 0 23.243562f
Cpar147 173 0 3.8650312f
Cpar148 174 0 3.24375f
Cpar149 175 0 3.3376875f
Cpar150 176 0 3.7905312f
Cpar151 177 0 3.6394063f
Cpar152 178 0 1.04175f
Cpar153 179 0 3.7905312f
Cpar154 180 0 3.24375f
Cpar155 181 0 3.2903437f
Cpar156 182 0 3.3376875f
Cpar157 185 0 2.52975f
Cpar158 186 0 4.0961875f
Cpar159 187 0 3.6394063f
Cpar160 188 0 23.243625f
Cpar161 189 0 3.8650312f
Cpar162 190 0 3.24375f
Cpar163 191 0 1.04175f
Cpar164 192 0 23.245625f
Cpar165 193 0 3.7905312f
Cpar166 194 0 2.52975f
Cpar167 195 0 4.0961875f
Cpar168 196 0 3.2903437f
Cpar169 197 0 3.3376875f
Cpar170 200 0 3.24375f
Cpar171 201 0 3.6394063f
Cpar172 202 0 3.8650312f
Cpar173 203 0 3.82275f
Cpar174 206 0 1.04175f
Cpar175 208 0 3.7905312f
Cpar176 209 0 2.52975f
Cpar177 210 0 4.0961875f
Cpar178 211 0 3.7905312f
Cpar179 212 0 2.52975f
Cpar180 213 0 4.0961875f
Cpar181 214 0 3.70775f
Cpar182 215 0 3.3040625f
Cpar183 216 0 3.2903437f
Cpar184 217 0 3.24375f
Cpar185 218 0 3.24375f
Cpar186 219 0 3.6394063f
Cpar187 220 0 23.351062f
Cpar188 221 0 12.786219f
Cpar189 222 0 22.174688f
Cpar190 224 0 3.2903437f
Cpar191 227 0 1.04175f
Cpar192 228 0 23.375438f
Cpar193 229 0 3.7905312f
Cpar194 230 0 2.52975f
Cpar195 231 0 4.0961875f
Cpar196 232 0 3.3911562f
Cpar197 233 0 3.24375f
Cpar198 234 0 3.6394063f
Cpar199 235 0 12.825703f
Cpar200 236 0 22.174688f
Cpar201 238 0 23.338394f
Cpar202 239 0 2.52975f
Cpar203 240 0 4.0961875f
Cpar204 241 0 3.7905312f
Cpar205 242 0 3.2859875f
Cpar206 243 0 3.24375f
Cpar207 244 0 3.3227344f
Cpar208 245 0 12.806188f
Cpar209 247 0 30.276625f
Cpar210 248 0 131.77105f
Cpar211 249 0 643.3195f
Cpar212 250 0 3.2903437f
Cpar213 251 0 3.82275f
Cpar214 252 0 3.3040625f
Cpar215 253 0 3.7905312f
Cpar216 256 0 1.04175f
Cpar217 257 0 4.0961875f
Cpar218 258 0 2.52975f
Cpar219 259 0 4.0961875f
Cpar220 260 0 3.7905312f
Cpar221 261 0 2.52975f
Cpar222 262 0 3.24375f
Cpar223 263 0 22.174688f
Cpar224 264 0 3.24375f
Cpar225 265 0 26.273344f
Cpar226 266 0 4.0961875f
Cpar227 267 0 3.7108438f
Cpar228 268 0 3.6394063f
Cpar229 269 0 12.786219f
Cpar230 271 0 1.04175f
Cpar231 272 0 3.82275f
Cpar232 273 0 3.2903437f
Cpar233 274 0 3.3040625f
Cpar234 275 0 3.7905312f
Cpar235 278 0 4.0961875f
Cpar236 279 0 2.52975f
Cpar237 280 0 4.0961875f
Cpar238 281 0 2.52975f
Cpar239 282 0 3.24375f
Cpar240 283 0 22.174688f
Cpar241 284 0 3.24375f
Cpar242 285 0 23.314469f
Cpar243 286 0 4.0961875f
Cpar244 288 0 3.7108438f
Cpar245 289 0 3.7905312f
Cpar246 290 0 12.786219f
Cpar247 291 0 3.82275f
Cpar248 292 0 3.6394063f
Cpar249 293 0 1.04175f
Cpar250 294 0 3.7905312f
Cpar251 295 0 3.7108438f
Cpar252 296 0 3.2903437f
Cpar253 297 0 3.3040625f
Cpar254 298 0 3.7905312f
Cpar255 301 0 4.0961875f
Cpar256 302 0 2.52975f
Cpar257 303 0 4.0961875f
Cpar258 304 0 2.52975f
Cpar259 305 0 3.6394063f
Cpar260 306 0 3.24375f
Cpar261 307 0 12.786219f
Cpar262 308 0 22.174688f
Cpar263 309 0 3.24375f
Cpar264 310 0 23.36075f
Cpar265 311 0 4.0961875f
Cpar266 313 0 3.82275f
Cpar267 314 0 1.04175f
Cpar268 315 0 4.0961875f
Cpar269 316 0 3.7905312f
Cpar270 317 0 2.52975f
Cpar271 318 0 4.0961875f
Cpar272 319 0 2.52975f
Cpar273 320 0 3.7108438f
Cpar274 321 0 3.2903437f
Cpar275 322 0 3.3040625f
Cpar276 323 0 4.0961875f
Cpar277 324 0 3.7905312f
Cpar278 327 0 3.24375f
Cpar279 328 0 3.6394063f
Cpar280 329 0 23.314469f
Cpar281 330 0 12.786219f
Cpar282 331 0 22.174688f
Cpar283 332 0 3.24375f
Cpar284 334 0 126.17797f
Cpar285 335 0 3.82275f
Cpar286 338 0 1.04175f
Cpar287 339 0 4.0961875f
Cpar288 340 0 3.7905312f
Cpar289 341 0 2.52975f
Cpar290 342 0 4.0961875f
Cpar291 343 0 2.52975f
Cpar292 344 0 3.7108438f
Cpar293 345 0 3.2903437f
Cpar294 346 0 3.3040625f
Cpar295 347 0 4.0961875f
Cpar296 348 0 3.7905312f
Cpar297 349 0 3.24375f
Cpar298 350 0 3.24375f
Cpar299 351 0 3.6394063f
Cpar300 352 0 12.786219f
Cpar301 353 0 22.174688f
Cpar302 354 0 23.365156f
Cpar303 356 0 3.2903437f
Cpar304 357 0 3.82275f
Cpar305 358 0 3.3040625f
Cpar306 361 0 1.04175f
Cpar307 362 0 4.0961875f
Cpar308 363 0 3.7905312f
Cpar309 364 0 2.52975f
Cpar310 365 0 4.0961875f
Cpar311 366 0 2.52975f
Cpar312 367 0 3.7108438f
Cpar313 368 0 3.24375f
Cpar314 369 0 3.24375f
Cpar315 370 0 4.0961875f
Cpar316 371 0 3.7905312f
Cpar317 372 0 3.6394063f
Cpar318 373 0 23.314469f
Cpar319 374 0 22.174688f
Cpar320 375 0 12.786219f
Cpar321 378 0 2.52975f
Cpar322 379 0 4.0961875f
Cpar323 380 0 3.7905312f
Cpar324 381 0 23.353831f
Cpar325 382 0 3.24375f
Cpar326 383 0 3.3302969f
Cpar327 384 0 12.806188f
Cpar328 386 0 643.3195f
Cpar329 387 0 74.2155f
Cpar330 388 0 3.2903437f
Cpar331 389 0 3.82275f
Cpar332 390 0 3.3040625f
Cpar333 393 0 1.04175f
Cpar334 394 0 4.0961875f
Cpar335 395 0 2.52975f
Cpar336 396 0 4.0961875f
Cpar337 397 0 3.7905312f
Cpar338 398 0 2.52975f
Cpar339 399 0 3.7905312f
Cpar340 400 0 3.24375f
Cpar341 401 0 3.24375f
Cpar342 402 0 22.174688f
Cpar343 403 0 27.053313f
Cpar344 404 0 3.732f
Cpar345 405 0 12.802406f
Cpar346 408 0 3.82275f
Cpar347 409 0 3.2903437f
Cpar348 410 0 3.3040625f
Cpar349 413 0 1.04175f
Cpar350 414 0 4.0961875f
Cpar351 415 0 2.52975f
Cpar352 416 0 4.0961875f
Cpar353 417 0 3.7905312f
Cpar354 418 0 2.52975f
Cpar355 419 0 3.7905312f
Cpar356 420 0 23.300875f
Cpar357 421 0 3.24375f
Cpar358 422 0 3.24375f
Cpar359 423 0 22.174688f
Cpar360 425 0 3.7316562f
Cpar361 427 0 23.288219f
Cpar362 428 0 12.802406f
Cpar363 429 0 12.786219f
Cpar364 430 0 3.82275f
Cpar365 431 0 1.04175f
Cpar366 432 0 3.7905312f
Cpar367 433 0 3.2903437f
Cpar368 434 0 3.3040625f
Cpar369 437 0 2.52975f
Cpar370 438 0 3.24375f
Cpar371 439 0 12.786219f
Cpar372 440 0 3.24375f
Cpar373 441 0 22.174688f
Cpar374 442 0 132.52867f
Cpar375 444 0 2.52975f
Cpar376 445 0 3.7316562f
Cpar377 447 0 4.0961875f
Cpar378 448 0 3.7905312f
Cpar379 449 0 4.0961875f
Cpar380 450 0 3.7905312f
Cpar381 451 0 12.802406f
Cpar382 452 0 3.82275f
Cpar383 453 0 1.04175f
Cpar384 454 0 3.7905312f
Cpar385 455 0 3.7905312f
Cpar386 456 0 2.52975f
Cpar387 457 0 3.7313125f
Cpar388 458 0 3.2903437f
Cpar389 459 0 3.3040625f
Cpar390 462 0 4.0961875f
Cpar391 463 0 3.24375f
Cpar392 464 0 2.52975f
Cpar393 465 0 4.0961875f
Cpar394 466 0 3.24375f
Cpar395 467 0 23.289531f
Cpar396 468 0 12.786219f
Cpar397 469 0 22.174688f
Cpar398 472 0 12.802406f
Cpar399 473 0 3.82275f
Cpar400 474 0 1.04175f
Cpar401 475 0 4.0961875f
Cpar402 476 0 3.7905312f
Cpar403 477 0 2.52975f
Cpar404 478 0 4.0961875f
Cpar405 479 0 3.7905312f
Cpar406 480 0 2.52975f
Cpar407 481 0 3.7316562f
Cpar408 482 0 3.2903437f
Cpar409 483 0 3.3040625f
Cpar410 486 0 3.24375f
Cpar411 487 0 3.24375f
Cpar412 488 0 12.786219f
Cpar413 489 0 22.174688f
Cpar414 490 0 23.333687f
Cpar415 493 0 12.802406f
Cpar416 494 0 3.82275f
Cpar417 495 0 3.3040625f
Cpar418 498 0 1.04175f
Cpar419 499 0 3.3040625f
Cpar420 500 0 4.0961875f
Cpar421 501 0 3.7905312f
Cpar422 502 0 3.2903437f
Cpar423 503 0 2.52975f
Cpar424 504 0 4.0961875f
Cpar425 505 0 3.7905312f
Cpar426 506 0 2.52975f
Cpar427 507 0 3.7316562f
Cpar428 508 0 3.24375f
Cpar429 509 0 3.24375f
Cpar430 510 0 12.802406f
Cpar431 511 0 23.289531f
Cpar432 512 0 12.786219f
Cpar433 515 0 3.7905312f
Cpar434 516 0 3.3322219f
Cpar435 518 0 2.52975f
Cpar436 519 0 4.0961875f
Cpar437 520 0 3.8650313f
Cpar438 521 0 22.980938f
Cpar439 522 0 23.326144f
Cpar440 523 0 3.24375f
Cpar441 524 0 12.825703f
Cpar442 526 0 74.2155f
Cpar443 527 0 20.365125f
Cpar444 528 0 3.3040625f
Cpar445 529 0 3.7905312f
Cpar446 530 0 3.82275f
Cpar447 532 0 2.52975f
Cpar448 533 0 2.52975f
Cpar449 534 0 4.0961875f
Cpar450 535 0 3.7905312f
Cpar451 536 0 27.554672f
Cpar452 537 0 28.980891f
Cpar453 538 0 3.24375f
Cpar454 539 0 22.174688f
Cpar455 540 0 3.24375f
Cpar456 541 0 3.6599375f
Cpar457 542 0 3.2903437f
Cpar458 543 0 3.3040625f
Cpar459 544 0 3.7905312f
Cpar460 545 0 3.82275f
Cpar461 548 0 1.04175f
Cpar462 549 0 4.0961875f
Cpar463 550 0 2.52975f
Cpar464 551 0 4.0961875f
Cpar465 552 0 3.7905312f
Cpar466 553 0 2.52975f
Cpar467 554 0 23.003313f
Cpar468 555 0 3.24375f
Cpar469 556 0 22.174688f
Cpar470 557 0 3.24375f
Cpar471 558 0 3.7275625f
Cpar472 559 0 4.4522813f
Cpar473 560 0 3.82275f
Cpar474 561 0 1.04175f
Cpar475 562 0 3.2903437f
Cpar476 563 0 3.3040625f
Cpar477 566 0 23.002f
Cpar478 567 0 3.24375f
Cpar479 568 0 4.975125f
Cpar480 569 0 22.174688f
Cpar481 570 0 2.52975f
Cpar482 571 0 3.24375f
Cpar483 572 0 2.52975f
Cpar484 573 0 3.7275625f
Cpar485 574 0 4.0961875f
Cpar486 575 0 3.7905312f
Cpar487 576 0 4.0961875f
Cpar488 577 0 3.82275f
Cpar489 578 0 1.04175f
Cpar490 579 0 3.7905312f
Cpar491 580 0 3.7275625f
Cpar492 581 0 3.3040625f
Cpar493 582 0 3.24375f
Cpar494 583 0 3.2903437f
Cpar495 584 0 3.7905312f
Cpar496 587 0 2.52975f
Cpar497 588 0 4.0961875f
Cpar498 589 0 3.24375f
Cpar499 590 0 2.52975f
Cpar500 591 0 4.0961875f
Cpar501 592 0 23.003313f
Cpar502 593 0 4.9761562f
Cpar503 594 0 22.174688f
Cpar504 595 0 3.82275f
Cpar505 596 0 1.04175f
Cpar506 597 0 2.52975f
Cpar507 598 0 4.0961875f
Cpar508 599 0 3.7905312f
Cpar509 600 0 2.52975f
Cpar510 601 0 4.0961875f
Cpar511 602 0 3.7279062f
Cpar512 603 0 3.3040625f
Cpar513 604 0 3.2903437f
Cpar514 605 0 3.24375f
Cpar515 606 0 3.7905312f
Cpar516 609 0 3.24375f
Cpar517 610 0 23.003313f
Cpar518 611 0 4.9761562f
Cpar519 612 0 22.174688f
Cpar520 613 0 3.82275f
Cpar521 616 0 1.04175f
Cpar522 617 0 2.52975f
Cpar523 618 0 3.3040625f
Cpar524 619 0 4.0961875f
Cpar525 620 0 3.7905312f
Cpar526 621 0 3.2903437f
Cpar527 622 0 2.52975f
Cpar528 623 0 4.0961875f
Cpar529 624 0 3.7279062f
Cpar530 625 0 3.24375f
Cpar531 626 0 3.7905312f
Cpar532 627 0 3.24375f
Cpar533 628 0 23.003313f
Cpar534 629 0 22.174688f
Cpar535 630 0 3.2903437f
Cpar536 633 0 1.04175f
Cpar537 634 0 4.0961875f
Cpar538 635 0 2.52975f
Cpar539 636 0 4.0961875f
Cpar540 637 0 3.7905312f
Cpar541 638 0 3.24375f
Cpar542 639 0 4.5894375f
Cpar543 640 0 44.412313f
Cpar544 641 0 20.365125f
Cpar545 642 0 30.276625f
Cpar546 643 0 44.412313f
Cpar547 644 0 120.49825f
Cpar548 645 0 3.82275f
Cpar549 646 0 3.3040625f
Cpar550 647 0 2.52975f
Cpar551 648 0 3.7905312f
Cpar552 649 0 3.24375f
Cpar553 650 0 22.174688f
Cpar554 651 0 3.82275f
Cpar555 652 0 3.3040625f
Cpar556 653 0 3.7905312f
Cpar557 654 0 3.24375f
Cpar558 655 0 22.174688f
Cpar559 656 0 2.52975f
Cpar560 657 0 3.82275f
Cpar561 658 0 3.7905312f
Cpar562 659 0 3.3040625f
Cpar563 660 0 3.24375f
Cpar564 661 0 2.52975f
Cpar565 662 0 22.174688f
Cpar566 663 0 3.82275f
Cpar567 664 0 3.7905312f
Cpar568 665 0 2.52975f
Cpar569 666 0 3.3040625f
Cpar570 667 0 3.24375f
Cpar571 668 0 22.174688f
Cpar572 669 0 3.82275f
Cpar573 670 0 3.7905312f
Cpar574 671 0 2.52975f
Cpar575 672 0 3.24375f
Cpar576 673 0 4.975125f
Cpar577 674 0 22.174688f
Cpar578 675 0 3.82275f
Cpar579 676 0 3.329875f
Cpar580 677 0 3.3040625f
Cpar581 678 0 2.52975f
Cpar582 679 0 3.7905312f
Cpar583 680 0 3.24375f
Cpar584 681 0 22.174688f
Cpar585 682 0 3.80175f
Cpar586 683 0 30.276625f
Cpar587 684 0 643.3195f
Cpar588 685 0 643.3195f
Cpar589 686 0 74.2155f
Cpar590 687 0 26.465641f
Cpar591 688 0 643.3195f
Cpar592 689 0 74.2155f
Cpar593 690 0 44.412313f
Cpar594 691 0 20.365125f
Cpar595 692 0 30.276625f
Cpar596 693 0 44.412313f
Cpar597 694 0 20.365125f
Cpar598 695 0 120.49825f
Cpar599 696 0 133.63656f
Cpar600 697 0 30.276625f
Cpar601 698 0 27.076828f
Cpar602 699 0 26.762125f
Cpar603 700 0 643.3195f
Cpar604 701 0 74.2155f
Cpar605 702 0 44.412313f
Cpar606 703 0 20.365125f
Cpar607 704 0 30.276625f
Cpar608 705 0 120.49825f
Cpar609 706 0 643.3195f
Cpar610 707 0 30.276625f
Cpar611 708 0 120.49825f
Cpar612 709 0 30.276625f
Cpar613 710 0 643.3195f
Cpar614 711 0 643.3195f
Cpar615 712 0 44.412313f
Cpar616 713 0 30.276625f
Cpar617 714 0 74.2155f
Cpar618 715 0 20.365125f
Cpar619 716 0 44.412313f
Cpar620 717 0 30.276625f
Cpar621 718 0 120.49825f
Cpar622 719 0 44.412313f
Cpar623 720 0 74.2155f
Cpar624 721 0 20.365125f
Cpar625 722 0 120.49825f
Cpar626 723 0 643.3195f
Cpar627 724 0 74.2155f
Cpar628 725 0 44.412312f
Cpar629 726 0 20.365125f
Cpar630 727 0 643.3195f
Cpar631 728 0 74.2155f
Cpar632 729 0 44.412313f
Cpar633 730 0 20.365125f
Cpar634 731 0 30.276625f
Cpar635 732 0 120.49825f
Cpar636 733 0 74.2155f
Cpar637 734 0 26.133406f
Cpar638 735 0 20.365125f
Cpar639 736 0 120.49825f
Cpar640 737 0 74.2155f
Cpar641 738 0 30.276625f
Cpar642 739 0 44.412312f
Cpar643 740 0 20.365125f
Cpar644 741 0 26.409781f
Cpar645 742 0 120.49825f
Cpar646 743 0 643.3195f
Cpar647 744 0 74.2155f
Cpar648 745 0 44.412313f
Cpar649 746 0 20.365125f
Cpar650 747 0 26.831047f
Cpar651 748 0 30.276625f
Cpar652 749 0 120.49825f
Cpar653 750 0 643.3195f

C4751 1 12  184.041f    ; (1133.5 788 1419.5 1074)CMOSN.041f    
C4747 2 12  184.041f    ; (697.5 788 983.5 1074)CMOSN.041f    
C4743 3 12  184.041f    ; (261.5 788 547.5 1074)CMOSN.041f    
C4739 4 12  184.041f    ; (-174.5 788 111.5 1074)CMOSN.041f    
C4735 5 12  184.041f    ; (-610.5 788 -324.5 1074)CMOSN.041f    
C4731 6 12  184.041f    ; (-1046.5 788 -760.5 1074)CMOSN.041f    
C4728 7 12  184.041f    ; (-1482.5 788 -1196.5 1074)CMOSN.041f    
M4725 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4724 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4723 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4722 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4721 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4720 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4719 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4718 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4717 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4716 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4715 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4714 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4712 are shorted:
* D4712 12 12 D_lateral AREA=3.249875f    ; (1408.5 613 1416.5 649)CMOSN4712 12 12 D_lateral AREA=3.249875f    
* Pins of element D4710 are shorted:
* D4710 12 12 D_lateral AREA=2.5E-016    ; (1392.5 648.999 1396.5 649)CMOSN4710 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4709 are shorted:
* D4709 12 12 D_lateral AREA=2.5E-016    ; (1376.5 648.999 1380.5 649)CMOSN4709 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4708 are shorted:
* D4708 12 12 D_lateral AREA=2.5E-016    ; (1360.5 648.999 1364.5 649)CMOSN4708 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4707 are shorted:
* D4707 12 12 D_lateral AREA=2.5E-016    ; (1344.5 648.999 1348.5 649)CMOSN4707 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4706 are shorted:
* D4706 12 12 D_lateral AREA=2.5E-016    ; (1328.5 648.999 1332.5 649)CMOSN4706 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4705 are shorted:
* D4705 12 12 D_lateral AREA=2.5E-016    ; (1312.5 648.999 1316.5 649)CMOSN4705 12 12 D_lateral AREA=2.5E-016    
M4702 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4701 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4700 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4699 1 11 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4689 are shorted:
* D4689 12 12 D_lateral AREA=2.5E-016    ; (1296.5 648.999 1300.5 649)CMOSN4689 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4688 are shorted:
* D4688 12 12 D_lateral AREA=2.3749375f    ; (1280.5 615 1284.5 649)CMOSN4688 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4677 are shorted:
* D4677 12 12 D_lateral AREA=2.5E-016    ; (1174.5 621.999 1178.5 622)CMOSN4677 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4676 are shorted:
* D4676 12 12 D_lateral AREA=2.5E-016    ; (1158.5 621.999 1162.5 622)CMOSN4676 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4675 are shorted:
* D4675 12 12 D_lateral AREA=2.5E-016    ; (1142.5 621.999 1146.5 622)CMOSN4675 12 12 D_lateral AREA=2.5E-016    
M4674 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4673 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4672 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4671 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4670 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4669 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4668 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4667 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4666 are shorted:
* D4666 12 12 D_lateral AREA=3.249875f    ; (972.5 613 980.5 649)CMOSN4666 12 12 D_lateral AREA=3.249875f    
* Pins of element D4665 are shorted:
* D4665 12 12 D_lateral AREA=2.5E-016    ; (956.5 648.999 960.5 649)CMOSN4665 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4664 are shorted:
* D4664 12 12 D_lateral AREA=2.5E-016    ; (940.5 648.999 944.5 649)CMOSN4664 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4663 are shorted:
* D4663 12 12 D_lateral AREA=2.5E-016    ; (924.5 648.999 928.5 649)CMOSN4663 12 12 D_lateral AREA=2.5E-016    
M4658 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4657 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4656 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4655 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4654 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4653 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4652 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4651 2 13 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4644 are shorted:
* D4644 12 12 D_lateral AREA=2.5E-016    ; (908.5 648.999 912.5 649)CMOSN4644 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4643 are shorted:
* D4643 12 12 D_lateral AREA=2.5E-016    ; (892.5 648.999 896.5 649)CMOSN4643 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4642 are shorted:
* D4642 12 12 D_lateral AREA=2.5E-016    ; (876.5 648.999 880.5 649)CMOSN4642 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4641 are shorted:
* D4641 12 12 D_lateral AREA=2.5E-016    ; (860.5 648.999 864.5 649)CMOSN4641 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4640 are shorted:
* D4640 12 12 D_lateral AREA=2.3749375f    ; (844.5 615 848.5 649)CMOSN4640 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4630 are shorted:
* D4630 12 12 D_lateral AREA=2f    ; (809.5 592.999 821.5 603)CMOSN4630 12 12 D_lateral AREA=2f    
* Pins of element D4626 are shorted:
* D4626 12 12 D_lateral AREA=2.5E-016    ; (738.5 621.999 742.5 622)CMOSN4626 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4625 are shorted:
* D4625 12 12 D_lateral AREA=2.5E-016    ; (722.5 621.999 726.5 622)CMOSN4625 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4623 are shorted:
* D4623 12 12 D_lateral AREA=2.5E-016    ; (706.5 621.999 710.5 622)CMOSN4623 12 12 D_lateral AREA=2.5E-016    
M4622 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4621 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4620 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4618 are shorted:
* D4618 12 12 D_lateral AREA=3.249875f    ; (536.5 613 544.5 649)CMOSN4618 12 12 D_lateral AREA=3.249875f    
* Pins of element D4617 are shorted:
* D4617 12 12 D_lateral AREA=2.5E-016    ; (520.5 648.999 524.5 649)CMOSN4617 12 12 D_lateral AREA=2.5E-016    
M4613 12 15 3 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4612 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4611 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4610 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4609 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4608 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4607 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4606 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4605 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4604 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4603 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4602 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4601 3 15 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4599 are shorted:
* D4599 12 12 D_lateral AREA=2.5E-016    ; (504.5 648.999 508.5 649)CMOSN4599 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4598 are shorted:
* D4598 12 12 D_lateral AREA=2.5E-016    ; (488.5 648.999 492.5 649)CMOSN4598 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4597 are shorted:
* D4597 12 12 D_lateral AREA=2.5E-016    ; (472.5 648.999 476.5 649)CMOSN4597 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4596 are shorted:
* D4596 12 12 D_lateral AREA=2.5E-016    ; (456.5 648.999 460.5 649)CMOSN4596 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4595 are shorted:
* D4595 12 12 D_lateral AREA=2.5E-016    ; (440.5 648.999 444.5 649)CMOSN4595 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4594 are shorted:
* D4594 12 12 D_lateral AREA=2.5E-016    ; (424.5 648.999 428.5 649)CMOSN4594 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4580 are shorted:
* D4580 12 12 D_lateral AREA=2.3749375f    ; (408.5 615 412.5 649)CMOSN4580 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4572 are shorted:
* D4572 12 12 D_lateral AREA=2.5E-016    ; (302.5 621.999 306.5 622)CMOSN4572 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4571 are shorted:
* D4571 12 12 D_lateral AREA=2.5E-016    ; (286.5 621.999 290.5 622)CMOSN4571 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4570 are shorted:
* D4570 12 12 D_lateral AREA=2.5E-016    ; (270.5 621.999 274.5 622)CMOSN4570 12 12 D_lateral AREA=2.5E-016    
M4569 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4568 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4567 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4566 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4565 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4564 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4563 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4562 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4561 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4560 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4559 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4557 are shorted:
* D4557 12 12 D_lateral AREA=3.249875f    ; (100.5 613 108.5 649)CMOSN4557 12 12 D_lateral AREA=3.249875f    
* Pins of element D4556 are shorted:
* D4556 12 12 D_lateral AREA=2.5E-016    ; (84.5 648.999 88.5 649)CMOSN4556 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4555 are shorted:
* D4555 12 12 D_lateral AREA=2.5E-016    ; (68.5 648.999 72.5 649)CMOSN4555 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4554 are shorted:
* D4554 12 12 D_lateral AREA=2.5E-016    ; (52.5 648.999 56.5 649)CMOSN4554 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4553 are shorted:
* D4553 12 12 D_lateral AREA=2.5E-016    ; (36.5 648.999 40.5 649)CMOSN4553 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4552 are shorted:
* D4552 12 12 D_lateral AREA=2.5E-016    ; (20.5 648.999 24.5 649)CMOSN4552 12 12 D_lateral AREA=2.5E-016    
M4548 12 21 4 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4547 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4546 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4545 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4544 4 21 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4535 are shorted:
* D4535 12 12 D_lateral AREA=2.5E-016    ; (4.5 648.999 8.5 649)CMOSN4535 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4534 are shorted:
* D4534 12 12 D_lateral AREA=2.5E-016    ; (-11.5 648.999 -7.5 649)CMOSN4534 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4533 are shorted:
* D4533 12 12 D_lateral AREA=2.3749375f    ; (-27.5 615 -23.5 649)CMOSN4533 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4521 are shorted:
* D4521 12 12 D_lateral AREA=2.5E-016    ; (-133.5 621.999 -129.5 622)CMOSN4521 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4520 are shorted:
* D4520 12 12 D_lateral AREA=2.5E-016    ; (-149.5 621.999 -145.5 622)CMOSN4520 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4519 are shorted:
* D4519 12 12 D_lateral AREA=2.5E-016    ; (-165.5 621.999 -161.5 622)CMOSN4519 12 12 D_lateral AREA=2.5E-016    
M4518 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4517 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4516 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4515 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4514 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4513 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4512 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4511 are shorted:
* D4511 12 12 D_lateral AREA=3.249875f    ; (-335.5 613 -327.5 649)CMOSN4511 12 12 D_lateral AREA=3.249875f    
* Pins of element D4510 are shorted:
* D4510 12 12 D_lateral AREA=2.5E-016    ; (-351.5 648.999 -347.5 649)CMOSN4510 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4509 are shorted:
* D4509 12 12 D_lateral AREA=2.5E-016    ; (-367.5 648.999 -363.5 649)CMOSN4509 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4508 are shorted:
* D4508 12 12 D_lateral AREA=2.5E-016    ; (-383.5 648.999 -379.5 649)CMOSN4508 12 12 D_lateral AREA=2.5E-016    
M4504 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4503 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4502 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4501 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4500 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4499 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4498 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4497 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4496 5 22 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4490 are shorted:
* D4490 12 12 D_lateral AREA=2.5E-016    ; (-399.5 648.999 -395.5 649)CMOSN4490 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4489 are shorted:
* D4489 12 12 D_lateral AREA=2.5E-016    ; (-415.5 648.999 -411.5 649)CMOSN4489 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4488 are shorted:
* D4488 12 12 D_lateral AREA=2.5E-016    ; (-431.5 648.999 -427.5 649)CMOSN4488 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4487 are shorted:
* D4487 12 12 D_lateral AREA=2.5E-016    ; (-447.5 648.999 -443.5 649)CMOSN4487 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4486 are shorted:
* D4486 12 12 D_lateral AREA=2.3749375f    ; (-463.5 615 -459.5 649)CMOSN4486 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4472 are shorted:
* D4472 12 12 D_lateral AREA=2.5E-016    ; (-569.5 621.999 -565.5 622)CMOSN4472 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4471 are shorted:
* D4471 12 12 D_lateral AREA=2.5E-016    ; (-585.5 621.999 -581.5 622)CMOSN4471 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4468 are shorted:
* D4468 12 12 D_lateral AREA=2.5E-016    ; (-601.5 621.999 -597.5 622)CMOSN4468 12 12 D_lateral AREA=2.5E-016    
M4467 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4466 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4464 are shorted:
* D4464 12 12 D_lateral AREA=3.249875f    ; (-771.5 613 -763.5 649)CMOSN4464 12 12 D_lateral AREA=3.249875f    
* Pins of element D4463 are shorted:
* D4463 12 12 D_lateral AREA=2.5E-016    ; (-787.5 648.999 -783.5 649)CMOSN4463 12 12 D_lateral AREA=2.5E-016    
M4459 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4458 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4457 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4456 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4455 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4454 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4453 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4452 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4451 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4450 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4449 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4448 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4447 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4446 are shorted:
* D4446 12 12 D_lateral AREA=2.5E-016    ; (-803.5 648.999 -799.5 649)CMOSN4446 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4445 are shorted:
* D4445 12 12 D_lateral AREA=2.5E-016    ; (-819.5 648.999 -815.5 649)CMOSN4445 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4444 are shorted:
* D4444 12 12 D_lateral AREA=2.5E-016    ; (-835.5 648.999 -831.5 649)CMOSN4444 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4443 are shorted:
* D4443 12 12 D_lateral AREA=2.5E-016    ; (-851.5 648.999 -847.5 649)CMOSN4443 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4442 are shorted:
* D4442 12 12 D_lateral AREA=2.5E-016    ; (-867.5 648.999 -863.5 649)CMOSN4442 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4441 are shorted:
* D4441 12 12 D_lateral AREA=2.5E-016    ; (-883.5 648.999 -879.5 649)CMOSN4441 12 12 D_lateral AREA=2.5E-016    
M4440 6 25 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4428 are shorted:
* D4428 12 12 D_lateral AREA=2.3749375f    ; (-899.5 615 -895.5 649)CMOSN4428 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4419 are shorted:
* D4419 12 12 D_lateral AREA=2.3749375f    ; (-989.5 588 -985.5 622)CMOSN4419 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4418 are shorted:
* D4418 12 12 D_lateral AREA=2.5E-016    ; (-1005.5 621.999 -1001.5 622)CMOSN4418 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4417 are shorted:
* D4417 12 12 D_lateral AREA=2.5E-016    ; (-1021.5 621.999 -1017.5 622)CMOSN4417 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4416 are shorted:
* D4416 12 12 D_lateral AREA=2.5E-016    ; (-1037.5 621.999 -1033.5 622)CMOSN4416 12 12 D_lateral AREA=2.5E-016    
M4415 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M4414 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4413 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4412 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4411 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4410 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4409 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4408 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4407 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4406 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D4404 are shorted:
* D4404 12 12 D_lateral AREA=3.249875f    ; (-1207.5 613 -1199.5 649)CMOSN4404 12 12 D_lateral AREA=3.249875f    
* Pins of element D4403 are shorted:
* D4403 12 12 D_lateral AREA=2.5E-016    ; (-1223.5 648.999 -1219.5 649)CMOSN4403 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4402 are shorted:
* D4402 12 12 D_lateral AREA=2.5E-016    ; (-1239.5 648.999 -1235.5 649)CMOSN4402 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4401 are shorted:
* D4401 12 12 D_lateral AREA=2.5E-016    ; (-1255.5 648.999 -1251.5 649)CMOSN4401 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4400 are shorted:
* D4400 12 12 D_lateral AREA=2.5E-016    ; (-1271.5 648.999 -1267.5 649)CMOSN4400 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4399 are shorted:
* D4399 12 12 D_lateral AREA=2.5E-016    ; (-1287.5 648.999 -1283.5 649)CMOSN4399 12 12 D_lateral AREA=2.5E-016    
M4395 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4394 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4393 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4392 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4391 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4390 7 30 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D4382 are shorted:
* D4382 12 12 D_lateral AREA=2.5E-016    ; (-1303.5 648.999 -1299.5 649)CMOSN4382 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4381 are shorted:
* D4381 12 12 D_lateral AREA=2.5E-016    ; (-1319.5 648.999 -1315.5 649)CMOSN4381 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4380 are shorted:
* D4380 12 12 D_lateral AREA=2.3749375f    ; (-1335.5 615 -1331.5 649)CMOSN4380 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4367 are shorted:
* D4367 12 12 D_lateral AREA=2.5E-016    ; (-1441.5 621.999 -1437.5 622)CMOSN4367 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4366 are shorted:
* D4366 12 12 D_lateral AREA=2.5E-016    ; (-1457.5 621.999 -1453.5 622)CMOSN4366 12 12 D_lateral AREA=2.5E-016    
* Pins of element D4365 are shorted:
* D4365 12 12 D_lateral AREA=2.5E-016    ; (-1473.5 621.999 -1469.5 622)CMOSN4365 12 12 D_lateral AREA=2.5E-016    
M4362 8 12 10 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M4360 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4358 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4356 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4354 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4352 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4350 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4348 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4346 1 10 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M4345 10 12 11 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
* Pins of element D4344 are shorted:
* D4344 8 8 D_lateral AREA=2.5E-016    ; (1395.5 589 1399.5 589.001)CMOSN4344 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4343 are shorted:
* D4343 8 8 D_lateral AREA=2.5E-016    ; (1379.5 589 1383.5 589.001)CMOSN4343 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4342 are shorted:
* D4342 8 8 D_lateral AREA=2.5E-016    ; (1363.5 589 1367.5 589.001)CMOSN4342 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4341 are shorted:
* D4341 8 8 D_lateral AREA=1.8125625f    ; (1345.499 566 1351.5 589.001)CMOSN4341 8 8 D_lateral AREA=1.8125625f    
* Pins of element D4340 are shorted:
* D4340 8 8 D_lateral AREA=3.5625625f    ; (1320.5 509.999 1330.501 557)CMOSN4340 8 8 D_lateral AREA=3.5625625f    
M4339 8 12 10 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M4338 8 12 10 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4337 10 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4336 31 1 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M4335 10 9 11 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M4334 11 9 10 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M4333 10 9 11 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M4332 9 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M4331 11 12 10 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M4330 10 12 11 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M4329 11 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M4328 11 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4327 12 12 11 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4326 11 9 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M4325 12 12 9 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
M4324 12 1 31 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
* Pins of element D4323 are shorted:
* D4323 12 12 D_lateral AREA=2f    ; (1245.5 592.999 1257.5 603)CMOSN4323 12 12 D_lateral AREA=2f    
* Pins of element D4322 are shorted:
* D4322 12 12 D_lateral AREA=3.75E-016    ; (1248.5 584 1254.5 584.001)CMOSN4322 12 12 D_lateral AREA=3.75E-016    
* Pins of element D4321 are shorted:
* D4321 12 12 D_lateral AREA=2.4374375f    ; (1214.5 586 1220.5 619)CMOSN4321 12 12 D_lateral AREA=2.4374375f    
* Pins of element D4320 are shorted:
* D4320 8 8 D_lateral AREA=4.1250625f    ; (1214.5 504 1222.501 562.001)CMOSN4320 8 8 D_lateral AREA=4.1250625f    
* Pins of element D4319 are shorted:
* D4319 8 8 D_lateral AREA=2.5E-016    ; (1304.5 509.999 1308.5 510)CMOSN4319 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4318 are shorted:
* D4318 8 8 D_lateral AREA=3.125E-016    ; (1287.5 509.999 1292.5 510)CMOSN4318 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4317 are shorted:
* D4317 8 8 D_lateral AREA=3.125E-016    ; (1287.5 563 1292.5 563.001)CMOSN4317 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4316 are shorted:
* D4316 8 8 D_lateral AREA=4.062625f    ; (1232.499 509.999 1238.5 563.001)CMOSN4316 8 8 D_lateral AREA=4.062625f    
M4315 8 31 73 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M4314 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4313 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4312 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4311 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4310 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4309 8 31 73 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M4308 31 1 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M4307 73 31 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M4306 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4305 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4304 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4303 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4302 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4301 12 31 73 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M4300 31 1 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D4299 are shorted:
* D4299 12 12 D_lateral AREA=2.687375f    ; (1198.5 586 1202.5 621)CMOSN4299 12 12 D_lateral AREA=2.687375f    
* Pins of element D4298 are shorted:
* D4298 12 12 D_lateral AREA=2.3749375f    ; (1190.5 588 1194.5 622)CMOSN4298 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4297 are shorted:
* D4297 8 8 D_lateral AREA=4.375E-016    ; (1194.5 562 1201.5 562.001)CMOSN4297 8 8 D_lateral AREA=4.375E-016    
M4294 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4292 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4290 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4288 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4286 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4284 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4282 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4280 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D4278 are shorted:
* D4278 8 8 D_lateral AREA=2.5E-016    ; (959.5 589 963.5 589.001)CMOSN4278 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4277 are shorted:
* D4277 8 8 D_lateral AREA=2.5E-016    ; (943.5 589 947.5 589.001)CMOSN4277 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4276 are shorted:
* D4276 8 8 D_lateral AREA=2.5E-016    ; (927.5 589 931.5 589.001)CMOSN4276 8 8 D_lateral AREA=2.5E-016    
M4274 32 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M4273 8 12 32 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4272 32 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4271 32 14 13 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M4270 13 14 32 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M4269 32 14 13 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M4268 8 12 32 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M4267 32 12 13 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M4266 13 12 32 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M4265 32 12 13 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M4264 13 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M4263 13 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4262 12 12 13 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4261 13 14 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D4259 are shorted:
* D4259 12 12 D_lateral AREA=3.75E-016    ; (812.5 584 818.5 584.001)CMOSN4259 12 12 D_lateral AREA=3.75E-016    
* Pins of element D4258 are shorted:
* D4258 8 8 D_lateral AREA=1.8125625f    ; (909.499 566 915.5 589.001)CMOSN4258 8 8 D_lateral AREA=1.8125625f    
* Pins of element D4257 are shorted:
* D4257 8 8 D_lateral AREA=3.5625625f    ; (884.5 509.999 894.501 557)CMOSN4257 8 8 D_lateral AREA=3.5625625f    
* Pins of element D4256 are shorted:
* D4256 8 8 D_lateral AREA=2.5E-016    ; (868.5 509.999 872.5 510)CMOSN4256 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4255 are shorted:
* D4255 8 8 D_lateral AREA=3.125E-016    ; (851.5 509.999 856.5 510)CMOSN4255 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4254 are shorted:
* D4254 8 8 D_lateral AREA=3.125E-016    ; (851.5 563 856.5 563.001)CMOSN4254 8 8 D_lateral AREA=3.125E-016    
M4253 8 33 83 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M4252 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4251 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4250 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4249 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4248 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4247 33 2 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M4246 33 2 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M4245 14 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M4244 83 33 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M4243 12 33 83 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4242 12 33 83 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4241 12 33 83 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4240 12 33 83 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4239 83 33 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M4238 12 12 14 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
M4237 33 2 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M4236 33 2 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D4235 are shorted:
* D4235 12 12 D_lateral AREA=2.4374375f    ; (778.5 586 784.5 619)CMOSN4235 12 12 D_lateral AREA=2.4374375f    
* Pins of element D4234 are shorted:
* D4234 12 12 D_lateral AREA=2.687375f    ; (762.5 586 766.5 621)CMOSN4234 12 12 D_lateral AREA=2.687375f    
* Pins of element D4233 are shorted:
* D4233 12 12 D_lateral AREA=2.3749375f    ; (754.5 588 758.5 622)CMOSN4233 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4232 are shorted:
* D4232 8 8 D_lateral AREA=4.1250625f    ; (778.5 504 786.501 562.001)CMOSN4232 8 8 D_lateral AREA=4.1250625f    
* Pins of element D4231 are shorted:
* D4231 8 8 D_lateral AREA=4.375E-016    ; (758.5 562 765.5 562.001)CMOSN4231 8 8 D_lateral AREA=4.375E-016    
* Pins of element D4229 are shorted:
* D4229 8 8 D_lateral AREA=4.062625f    ; (796.499 509.999 802.5 563.001)CMOSN4229 8 8 D_lateral AREA=4.062625f    
M4228 8 33 83 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M4227 12 33 83 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M4225 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4223 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4221 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4219 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D4217 are shorted:
* D4217 8 8 D_lateral AREA=2.5E-016    ; (523.5 589 527.5 589.001)CMOSN4217 8 8 D_lateral AREA=2.5E-016    
M4215 34 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M4214 8 12 34 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4213 34 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4212 8 12 34 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M4210 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4208 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4206 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4204 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M4203 34 12 15 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M4202 15 12 34 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M4201 34 12 15 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
* Pins of element D4199 are shorted:
* D4199 8 8 D_lateral AREA=2.5E-016    ; (507.5 589 511.5 589.001)CMOSN4199 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4198 are shorted:
* D4198 8 8 D_lateral AREA=2.5E-016    ; (491.5 589 495.5 589.001)CMOSN4198 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4197 are shorted:
* D4197 8 8 D_lateral AREA=1.8125625f    ; (473.499 566 479.5 589.001)CMOSN4197 8 8 D_lateral AREA=1.8125625f    
* Pins of element D4196 are shorted:
* D4196 8 8 D_lateral AREA=3.5625625f    ; (448.5 509.999 458.501 557)CMOSN4196 8 8 D_lateral AREA=3.5625625f    
* Pins of element D4195 are shorted:
* D4195 8 8 D_lateral AREA=2.5E-016    ; (432.5 509.999 436.5 510)CMOSN4195 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4194 are shorted:
* D4194 8 8 D_lateral AREA=3.125E-016    ; (415.5 509.999 420.5 510)CMOSN4194 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4193 are shorted:
* D4193 8 8 D_lateral AREA=3.125E-016    ; (415.5 563 420.5 563.001)CMOSN4193 8 8 D_lateral AREA=3.125E-016    
M4192 8 17 18 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M4191 17 3 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M4190 17 3 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M4189 34 16 15 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M4188 15 16 34 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M4187 34 16 15 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M4186 16 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M4185 12 17 18 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M4184 15 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M4183 15 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4182 12 12 15 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4181 15 16 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M4180 12 12 16 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
M4179 17 3 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M4178 17 3 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D4177 are shorted:
* D4177 12 12 D_lateral AREA=2f    ; (373.5 592.999 385.5 603)CMOSN4177 12 12 D_lateral AREA=2f    
* Pins of element D4176 are shorted:
* D4176 12 12 D_lateral AREA=3.75E-016    ; (376.5 584 382.5 584.001)CMOSN4176 12 12 D_lateral AREA=3.75E-016    
* Pins of element D4175 are shorted:
* D4175 12 12 D_lateral AREA=2.4374375f    ; (342.5 586 348.5 619)CMOSN4175 12 12 D_lateral AREA=2.4374375f    
* Pins of element D4174 are shorted:
* D4174 12 12 D_lateral AREA=2.687375f    ; (326.5 586 330.5 621)CMOSN4174 12 12 D_lateral AREA=2.687375f    
* Pins of element D4173 are shorted:
* D4173 12 12 D_lateral AREA=2.3749375f    ; (318.5 588 322.5 622)CMOSN4173 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4172 are shorted:
* D4172 8 8 D_lateral AREA=4.1250625f    ; (342.5 504 350.501 562.001)CMOSN4172 8 8 D_lateral AREA=4.1250625f    
* Pins of element D4171 are shorted:
* D4171 8 8 D_lateral AREA=4.375E-016    ; (322.5 562 329.5 562.001)CMOSN4171 8 8 D_lateral AREA=4.375E-016    
* Pins of element D4169 are shorted:
* D4169 8 8 D_lateral AREA=4.062625f    ; (360.499 509.999 366.5 563.001)CMOSN4169 8 8 D_lateral AREA=4.062625f    
M4168 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4167 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4166 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4165 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4164 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4163 8 17 18 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M4162 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4161 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4160 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4159 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4158 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4157 12 17 18 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M4154 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4152 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4150 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4148 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4146 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4144 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4142 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4140 4 20 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D4138 are shorted:
* D4138 8 8 D_lateral AREA=2.5E-016    ; (87.5 589 91.5 589.001)CMOSN4138 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4137 are shorted:
* D4137 8 8 D_lateral AREA=2.5E-016    ; (71.5 589 75.5 589.001)CMOSN4137 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4136 are shorted:
* D4136 8 8 D_lateral AREA=2.5E-016    ; (55.5 589 59.5 589.001)CMOSN4136 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4135 are shorted:
* D4135 8 8 D_lateral AREA=1.8125625f    ; (37.499 566 43.5 589.001)CMOSN4135 8 8 D_lateral AREA=1.8125625f    
* Pins of element D4134 are shorted:
* D4134 8 8 D_lateral AREA=3.5625625f    ; (12.5 509.999 22.501 557)CMOSN4134 8 8 D_lateral AREA=3.5625625f    
M4133 20 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M4132 8 12 20 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4131 20 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4130 20 19 21 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M4129 21 19 20 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M4128 20 19 21 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M4127 19 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M4126 20 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M4125 20 12 21 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M4124 21 12 20 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M4123 20 12 21 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M4122 21 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M4121 21 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4120 12 12 21 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4119 21 19 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M4118 12 12 19 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
* Pins of element D4117 are shorted:
* D4117 12 12 D_lateral AREA=2f    ; (-62.5 592.999 -50.5 603)CMOSN4117 12 12 D_lateral AREA=2f    
* Pins of element D4116 are shorted:
* D4116 12 12 D_lateral AREA=3.75E-016    ; (-59.5 584 -53.5 584.001)CMOSN4116 12 12 D_lateral AREA=3.75E-016    
* Pins of element D4113 are shorted:
* D4113 8 8 D_lateral AREA=2.5E-016    ; (-3.5 509.999 0.5 510)CMOSN4113 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4112 are shorted:
* D4112 8 8 D_lateral AREA=3.125E-016    ; (-20.5 509.999 -15.5 510)CMOSN4112 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4111 are shorted:
* D4111 8 8 D_lateral AREA=3.125E-016    ; (-20.5 563 -15.5 563.001)CMOSN4111 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4110 are shorted:
* D4110 8 8 D_lateral AREA=4.062625f    ; (-75.501 509.999 -69.5 563.001)CMOSN4110 8 8 D_lateral AREA=4.062625f    
M4109 8 35 334 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M4108 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4107 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4106 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4105 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4104 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4103 8 35 334 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M4102 35 4 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M4101 35 4 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M4100 334 35 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M4099 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4098 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4097 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4096 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4095 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4094 12 35 334 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M4093 35 4 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M4092 35 4 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D4091 are shorted:
* D4091 12 12 D_lateral AREA=2.4374375f    ; (-93.5 586 -87.5 619)CMOSN4091 12 12 D_lateral AREA=2.4374375f    
* Pins of element D4090 are shorted:
* D4090 12 12 D_lateral AREA=2.687375f    ; (-109.5 586 -105.5 621)CMOSN4090 12 12 D_lateral AREA=2.687375f    
* Pins of element D4089 are shorted:
* D4089 12 12 D_lateral AREA=2.3749375f    ; (-117.5 588 -113.5 622)CMOSN4089 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4088 are shorted:
* D4088 8 8 D_lateral AREA=4.1250625f    ; (-93.5 504 -85.499 562.001)CMOSN4088 8 8 D_lateral AREA=4.1250625f    
* Pins of element D4087 are shorted:
* D4087 8 8 D_lateral AREA=4.375E-016    ; (-113.5 562 -106.5 562.001)CMOSN4087 8 8 D_lateral AREA=4.375E-016    
M4084 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4082 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4080 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4078 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4076 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4074 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4072 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D4070 are shorted:
* D4070 8 8 D_lateral AREA=2.5E-016    ; (-348.5 589 -344.5 589.001)CMOSN4070 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4069 are shorted:
* D4069 8 8 D_lateral AREA=2.5E-016    ; (-364.5 589 -360.5 589.001)CMOSN4069 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4068 are shorted:
* D4068 8 8 D_lateral AREA=2.5E-016    ; (-380.5 589 -376.5 589.001)CMOSN4068 8 8 D_lateral AREA=2.5E-016    
M4067 36 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M4066 8 12 36 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4065 36 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4064 36 23 22 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M4063 22 23 36 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M4062 36 23 22 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M4061 8 12 36 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M4059 5 36 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M4058 36 12 22 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M4057 22 12 36 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M4056 36 12 22 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M4055 22 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M4054 22 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4053 12 12 22 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M4052 22 23 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D4051 are shorted:
* D4051 8 8 D_lateral AREA=1.8125625f    ; (-398.501 566 -392.5 589.001)CMOSN4051 8 8 D_lateral AREA=1.8125625f    
* Pins of element D4050 are shorted:
* D4050 8 8 D_lateral AREA=3.5625625f    ; (-423.5 509.999 -413.499 557)CMOSN4050 8 8 D_lateral AREA=3.5625625f    
* Pins of element D4049 are shorted:
* D4049 8 8 D_lateral AREA=2.5E-016    ; (-439.5 509.999 -435.5 510)CMOSN4049 8 8 D_lateral AREA=2.5E-016    
* Pins of element D4048 are shorted:
* D4048 8 8 D_lateral AREA=3.125E-016    ; (-456.5 509.999 -451.5 510)CMOSN4048 8 8 D_lateral AREA=3.125E-016    
* Pins of element D4047 are shorted:
* D4047 8 8 D_lateral AREA=3.125E-016    ; (-456.5 563 -451.5 563.001)CMOSN4047 8 8 D_lateral AREA=3.125E-016    
M4046 8 24 37 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M4045 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4044 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4043 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4042 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4041 24 5 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M4040 24 5 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M4039 23 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M4038 37 24 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M4037 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4036 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4035 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4034 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4033 12 12 23 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
M4032 24 5 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M4031 24 5 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D4030 are shorted:
* D4030 12 12 D_lateral AREA=2f    ; (-498.5 592.999 -486.5 603)CMOSN4030 12 12 D_lateral AREA=2f    
* Pins of element D4029 are shorted:
* D4029 12 12 D_lateral AREA=3.75E-016    ; (-495.5 584 -489.5 584.001)CMOSN4029 12 12 D_lateral AREA=3.75E-016    
* Pins of element D4028 are shorted:
* D4028 12 12 D_lateral AREA=2.4374375f    ; (-529.5 586 -523.5 619)CMOSN4028 12 12 D_lateral AREA=2.4374375f    
* Pins of element D4027 are shorted:
* D4027 12 12 D_lateral AREA=2.687375f    ; (-545.5 586 -541.5 621)CMOSN4027 12 12 D_lateral AREA=2.687375f    
* Pins of element D4026 are shorted:
* D4026 12 12 D_lateral AREA=2.3749375f    ; (-553.5 588 -549.5 622)CMOSN4026 12 12 D_lateral AREA=2.3749375f    
* Pins of element D4025 are shorted:
* D4025 8 8 D_lateral AREA=4.1250625f    ; (-529.5 504 -521.499 562.001)CMOSN4025 8 8 D_lateral AREA=4.1250625f    
* Pins of element D4024 are shorted:
* D4024 8 8 D_lateral AREA=4.375E-016    ; (-549.5 562 -542.5 562.001)CMOSN4024 8 8 D_lateral AREA=4.375E-016    
* Pins of element D4022 are shorted:
* D4022 8 8 D_lateral AREA=4.062625f    ; (-511.501 509.999 -505.5 563.001)CMOSN4022 8 8 D_lateral AREA=4.062625f    
M4021 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M4020 8 24 37 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M4019 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M4018 12 24 37 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M4016 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M4014 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4012 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D4010 are shorted:
* D4010 8 8 D_lateral AREA=2.5E-016    ; (-784.5 589 -780.5 589.001)CMOSN4010 8 8 D_lateral AREA=2.5E-016    
M4009 27 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M4008 8 12 27 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M4007 27 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M4006 8 12 27 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M4004 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4002 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M4000 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3998 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3996 6 27 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M3995 27 12 25 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M3994 25 12 27 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M3993 27 12 25 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
* Pins of element D3992 are shorted:
* D3992 8 8 D_lateral AREA=2.5E-016    ; (-800.5 589 -796.5 589.001)CMOSN3992 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3991 are shorted:
* D3991 8 8 D_lateral AREA=2.5E-016    ; (-816.5 589 -812.5 589.001)CMOSN3991 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3990 are shorted:
* D3990 8 8 D_lateral AREA=1.8125625f    ; (-834.501 566 -828.5 589.001)CMOSN3990 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3989 are shorted:
* D3989 8 8 D_lateral AREA=3.5625625f    ; (-859.5 509.999 -849.499 557)CMOSN3989 8 8 D_lateral AREA=3.5625625f    
* Pins of element D3988 are shorted:
* D3988 8 8 D_lateral AREA=2.5E-016    ; (-875.5 509.999 -871.5 510)CMOSN3988 8 8 D_lateral AREA=2.5E-016    
M3985 38 6 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M3984 38 6 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3983 27 26 25 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M3982 25 26 27 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3981 27 26 25 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M3980 26 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M3979 25 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M3978 25 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3977 12 12 25 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3976 25 26 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M3975 12 12 26 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
M3974 38 6 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M3973 38 6 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D3972 are shorted:
* D3972 12 12 D_lateral AREA=2f    ; (-934.5 592.999 -922.5 603)CMOSN3972 12 12 D_lateral AREA=2f    
* Pins of element D3971 are shorted:
* D3971 12 12 D_lateral AREA=3.75E-016    ; (-931.5 584 -925.5 584.001)CMOSN3971 12 12 D_lateral AREA=3.75E-016    
* Pins of element D3970 are shorted:
* D3970 12 12 D_lateral AREA=2.4374375f    ; (-965.5 586 -959.5 619)CMOSN3970 12 12 D_lateral AREA=2.4374375f    
* Pins of element D3969 are shorted:
* D3969 12 12 D_lateral AREA=2.687375f    ; (-981.5 586 -977.5 621)CMOSN3969 12 12 D_lateral AREA=2.687375f    
* Pins of element D3967 are shorted:
* D3967 8 8 D_lateral AREA=4.1250625f    ; (-965.5 504 -957.499 562.001)CMOSN3967 8 8 D_lateral AREA=4.1250625f    
* Pins of element D3966 are shorted:
* D3966 8 8 D_lateral AREA=4.375E-016    ; (-985.5 562 -978.5 562.001)CMOSN3966 8 8 D_lateral AREA=4.375E-016    
* Pins of element D3964 are shorted:
* D3964 8 8 D_lateral AREA=3.125E-016    ; (-892.5 509.999 -887.5 510)CMOSN3964 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3963 are shorted:
* D3963 8 8 D_lateral AREA=3.125E-016    ; (-892.5 563 -887.5 563.001)CMOSN3963 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3962 are shorted:
* D3962 8 8 D_lateral AREA=4.062625f    ; (-947.501 509.999 -941.5 563.001)CMOSN3962 8 8 D_lateral AREA=4.062625f    
M3961 8 38 40 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M3960 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3959 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3958 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3957 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3956 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3955 8 38 40 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M3954 12 38 40 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M3953 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3952 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3951 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3950 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3949 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3948 12 38 40 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M3946 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3944 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3942 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3940 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3938 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3936 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3934 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3932 7 29 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D3930 are shorted:
* D3930 8 8 D_lateral AREA=2.5E-016    ; (-1220.5 589 -1216.5 589.001)CMOSN3930 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3929 are shorted:
* D3929 8 8 D_lateral AREA=2.5E-016    ; (-1236.5 589 -1232.5 589.001)CMOSN3929 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3928 are shorted:
* D3928 8 8 D_lateral AREA=2.5E-016    ; (-1252.5 589 -1248.5 589.001)CMOSN3928 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3927 are shorted:
* D3927 8 8 D_lateral AREA=1.8125625f    ; (-1270.501 566 -1264.5 589.001)CMOSN3927 8 8 D_lateral AREA=1.8125625f    
M3925 29 12 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M3924 8 12 29 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M3923 29 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M3922 29 28 30 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M3921 30 28 29 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3920 29 28 30 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M3919 28 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M3918 8 12 29 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M3917 29 12 30 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M3916 30 12 29 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M3915 29 12 30 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M3914 30 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M3913 30 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3912 12 12 30 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3911 30 28 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M3910 12 12 28 12 CMOSN L=500n W=3.75u AD=6.0625p PD=10.75u AS=5.625p PS=10.5u    
* Pins of element D3909 are shorted:
* D3909 12 12 D_lateral AREA=2f    ; (-1370.5 592.999 -1358.5 603)CMOSN3909 12 12 D_lateral AREA=2f    
* Pins of element D3908 are shorted:
* D3908 12 12 D_lateral AREA=3.75E-016    ; (-1367.5 584 -1361.5 584.001)CMOSN3908 12 12 D_lateral AREA=3.75E-016    
* Pins of element D3907 are shorted:
* D3907 8 8 D_lateral AREA=3.5625625f    ; (-1295.5 509.999 -1285.499 557)CMOSN3907 8 8 D_lateral AREA=3.5625625f    
* Pins of element D3906 are shorted:
* D3906 8 8 D_lateral AREA=2.5E-016    ; (-1311.5 509.999 -1307.5 510)CMOSN3906 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3905 are shorted:
* D3905 8 8 D_lateral AREA=3.125E-016    ; (-1328.5 509.999 -1323.5 510)CMOSN3905 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3904 are shorted:
* D3904 8 8 D_lateral AREA=3.125E-016    ; (-1328.5 563 -1323.5 563.001)CMOSN3904 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3903 are shorted:
* D3903 8 8 D_lateral AREA=4.062625f    ; (-1383.501 509.999 -1377.5 563.001)CMOSN3903 8 8 D_lateral AREA=4.062625f    
M3902 8 39 41 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M3901 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3900 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3899 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3898 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3897 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3896 8 39 41 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M3895 39 7 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M3894 39 7 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3893 41 39 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3892 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3891 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3890 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3889 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3888 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3887 12 39 41 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M3886 39 7 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M3885 39 7 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D3884 are shorted:
* D3884 12 12 D_lateral AREA=2.4374375f    ; (-1401.5 586 -1395.5 619)CMOSN3884 12 12 D_lateral AREA=2.4374375f    
* Pins of element D3883 are shorted:
* D3883 12 12 D_lateral AREA=2.687375f    ; (-1417.5 586 -1413.5 621)CMOSN3883 12 12 D_lateral AREA=2.687375f    
* Pins of element D3882 are shorted:
* D3882 12 12 D_lateral AREA=2.3749375f    ; (-1425.5 588 -1421.5 622)CMOSN3882 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3881 are shorted:
* D3881 8 8 D_lateral AREA=4.1250625f    ; (-1401.5 504 -1393.499 562.001)CMOSN3881 8 8 D_lateral AREA=4.1250625f    
* Pins of element D3880 are shorted:
* D3880 8 8 D_lateral AREA=4.375E-016    ; (-1421.5 562 -1414.5 562.001)CMOSN3880 8 8 D_lateral AREA=4.375E-016    
* Pins of element D3878 are shorted:
* D3878 8 8 D_lateral AREA=8.875125f    ; (1411.5 453.999 1415.501 589.001)CMOSN3878 8 8 D_lateral AREA=8.875125f    
M3877 8 10 1 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3876 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3875 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3874 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3873 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3872 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3871 8 10 1 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3870 8 10 1 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3869 are shorted:
* D3869 8 8 D_lateral AREA=8.625f    ; (1190.5 493.999 1202.5 557)CMOSN3869 8 8 D_lateral AREA=8.625f    
* Pins of element D3867 are shorted:
* D3867 8 8 D_lateral AREA=2.5E-016    ; (1174.5 493.999 1178.5 494)CMOSN3867 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3866 are shorted:
* D3866 8 8 D_lateral AREA=2.5E-016    ; (1158.5 493.999 1162.5 494)CMOSN3866 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3865 are shorted:
* D3865 8 8 D_lateral AREA=2.5E-016    ; (1142.5 493.999 1146.5 494)CMOSN3865 8 8 D_lateral AREA=2.5E-016    
M3864 8 32 2 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3863 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3862 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3861 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3860 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3859 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3858 8 32 2 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3857 2 32 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D3856 are shorted:
* D3856 8 8 D_lateral AREA=8.875125f    ; (975.5 453.999 979.501 589.001)CMOSN3856 8 8 D_lateral AREA=8.875125f    
* Pins of element D3855 are shorted:
* D3855 8 8 D_lateral AREA=8.625f    ; (754.5 493.999 766.5 557)CMOSN3855 8 8 D_lateral AREA=8.625f    
* Pins of element D3853 are shorted:
* D3853 8 8 D_lateral AREA=2.5E-016    ; (738.5 493.999 742.5 494)CMOSN3853 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3852 are shorted:
* D3852 8 8 D_lateral AREA=2.5E-016    ; (722.5 493.999 726.5 494)CMOSN3852 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3851 are shorted:
* D3851 8 8 D_lateral AREA=2.5E-016    ; (706.5 493.999 710.5 494)CMOSN3851 8 8 D_lateral AREA=2.5E-016    
M3850 8 34 3 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3849 8 34 3 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3848 8 34 3 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3847 3 34 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D3846 are shorted:
* D3846 8 8 D_lateral AREA=8.875125f    ; (539.5 453.999 543.501 589.001)CMOSN3846 8 8 D_lateral AREA=8.875125f    
M3845 8 34 3 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3844 8 34 3 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3843 8 34 3 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3842 8 34 3 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3841 are shorted:
* D3841 8 8 D_lateral AREA=8.625f    ; (318.5 493.999 330.5 557)CMOSN3841 8 8 D_lateral AREA=8.625f    
* Pins of element D3839 are shorted:
* D3839 8 8 D_lateral AREA=2.5E-016    ; (302.5 493.999 306.5 494)CMOSN3839 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3838 are shorted:
* D3838 8 8 D_lateral AREA=2.5E-016    ; (286.5 493.999 290.5 494)CMOSN3838 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3837 are shorted:
* D3837 8 8 D_lateral AREA=2.5E-016    ; (270.5 493.999 274.5 494)CMOSN3837 8 8 D_lateral AREA=2.5E-016    
M3836 8 20 4 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3835 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3834 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3833 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3832 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3831 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3830 8 20 4 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3829 8 20 4 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3828 are shorted:
* D3828 8 8 D_lateral AREA=8.875125f    ; (103.5 453.999 107.501 589.001)CMOSN3828 8 8 D_lateral AREA=8.875125f    
* Pins of element D3827 are shorted:
* D3827 8 8 D_lateral AREA=8.625f    ; (-117.5 493.999 -105.5 557)CMOSN3827 8 8 D_lateral AREA=8.625f    
* Pins of element D3825 are shorted:
* D3825 8 8 D_lateral AREA=2.5E-016    ; (-133.5 493.999 -129.5 494)CMOSN3825 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3824 are shorted:
* D3824 8 8 D_lateral AREA=2.5E-016    ; (-149.5 493.999 -145.5 494)CMOSN3824 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3823 are shorted:
* D3823 8 8 D_lateral AREA=2.5E-016    ; (-165.5 493.999 -161.5 494)CMOSN3823 8 8 D_lateral AREA=2.5E-016    
M3822 8 36 5 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3821 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3820 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3819 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3818 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3817 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3816 8 36 5 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D3815 are shorted:
* D3815 8 8 D_lateral AREA=8.875125f    ; (-332.5 453.999 -328.499 589.001)CMOSN3815 8 8 D_lateral AREA=8.875125f    
M3814 8 36 5 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3813 are shorted:
* D3813 8 8 D_lateral AREA=8.625f    ; (-553.5 493.999 -541.5 557)CMOSN3813 8 8 D_lateral AREA=8.625f    
* Pins of element D3811 are shorted:
* D3811 8 8 D_lateral AREA=2.5E-016    ; (-569.5 493.999 -565.5 494)CMOSN3811 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3810 are shorted:
* D3810 8 8 D_lateral AREA=2.5E-016    ; (-585.5 493.999 -581.5 494)CMOSN3810 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3809 are shorted:
* D3809 8 8 D_lateral AREA=2.5E-016    ; (-601.5 493.999 -597.5 494)CMOSN3809 8 8 D_lateral AREA=2.5E-016    
M3808 8 27 6 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3807 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3806 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D3805 are shorted:
* D3805 8 8 D_lateral AREA=8.875125f    ; (-768.5 453.999 -764.499 589.001)CMOSN3805 8 8 D_lateral AREA=8.875125f    
M3804 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3803 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3802 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3801 8 27 6 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3800 8 27 6 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3799 are shorted:
* D3799 8 8 D_lateral AREA=8.625f    ; (-989.5 493.999 -977.5 557)CMOSN3799 8 8 D_lateral AREA=8.625f    
* Pins of element D3796 are shorted:
* D3796 8 8 D_lateral AREA=2.5E-016    ; (-1005.5 493.999 -1001.5 494)CMOSN3796 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3795 are shorted:
* D3795 8 8 D_lateral AREA=2.5E-016    ; (-1021.5 493.999 -1017.5 494)CMOSN3795 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3794 are shorted:
* D3794 8 8 D_lateral AREA=2.5E-016    ; (-1037.5 493.999 -1033.5 494)CMOSN3794 8 8 D_lateral AREA=2.5E-016    
M3793 8 29 7 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M3792 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3791 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3790 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3789 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3788 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3787 8 29 7 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3786 8 29 7 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D3785 are shorted:
* D3785 8 8 D_lateral AREA=8.875125f    ; (-1204.5 453.999 -1200.499 589.001)CMOSN3785 8 8 D_lateral AREA=8.875125f    
* Pins of element D3784 are shorted:
* D3784 8 8 D_lateral AREA=8.625f    ; (-1425.5 493.999 -1413.5 557)CMOSN3784 8 8 D_lateral AREA=8.625f    
* Pins of element D3782 are shorted:
* D3782 8 8 D_lateral AREA=2.5E-016    ; (-1441.5 493.999 -1437.5 494)CMOSN3782 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3781 are shorted:
* D3781 8 8 D_lateral AREA=2.5E-016    ; (-1457.5 493.999 -1453.5 494)CMOSN3781 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3780 are shorted:
* D3780 8 8 D_lateral AREA=2.5E-016    ; (-1473.5 493.999 -1469.5 494)CMOSN3780 8 8 D_lateral AREA=2.5E-016    
M3766 8 42 47 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3764 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3762 8 42 47 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3760 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3758 8 42 47 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3756 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3754 8 42 47 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3752 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3748 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M3747 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3746 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3745 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3744 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3743 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3742 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3741 47 42 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3739 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3738 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3737 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3736 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3735 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3734 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3733 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3732 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D3731 are shorted:
* D3731 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 296 -1760.499 300)CMOSN3731 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3730 are shorted:
* D3730 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 312 -1760.499 316)CMOSN3730 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3729 are shorted:
* D3729 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 328 -1760.499 332)CMOSN3729 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3728 are shorted:
* D3728 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 344 -1760.499 348)CMOSN3728 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3727 are shorted:
* D3727 12 12 D_lateral AREA=3.249875f    ; (-1760.5 360 -1724.5 368)CMOSN3727 12 12 D_lateral AREA=3.249875f    
* Pins of element D3726 are shorted:
* D3726 8 8 D_lateral AREA=1.8125625f    ; (-1700.501 296.999 -1677.5 303)CMOSN3726 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3725 are shorted:
* D3725 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 315 -1700.5 319)CMOSN3725 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3724 are shorted:
* D3724 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 331 -1700.5 335)CMOSN3724 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3723 are shorted:
* D3723 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 347 -1700.5 351)CMOSN3723 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3722 are shorted:
* D3722 8 8 D_lateral AREA=8.875125f    ; (-1700.501 363 -1565.499 367.001)CMOSN3722 8 8 D_lateral AREA=8.875125f    
M3714 8 12 42 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M3713 42 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M3712 42 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M3711 43 44 42 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M3710 42 44 43 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3709 43 44 42 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M3708 42 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
* Pins of element D3707 are shorted:
* D3707 8 8 D_lateral AREA=2.5E-016    ; (-1621.5 256 -1621.499 260)CMOSN3707 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3706 are shorted:
* D3706 8 8 D_lateral AREA=3.5625625f    ; (-1668.5 272 -1621.499 282.001)CMOSN3706 8 8 D_lateral AREA=3.5625625f    
* Pins of element D3705 are shorted:
* D3705 8 8 D_lateral AREA=3.125E-016    ; (-1621.5 239 -1621.499 244)CMOSN3705 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3704 are shorted:
* D3704 8 8 D_lateral AREA=3.125E-016    ; (-1674.501 239 -1674.5 244)CMOSN3704 8 8 D_lateral AREA=3.125E-016    
M3703 43 12 42 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M3702 42 12 43 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M3701 43 12 42 12 CMOSN L=500n W=3.25u AD=2.53125p PD=5u AS=4.875p PS=9.5u    
M3700 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3699 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3698 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3697 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3696 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3695 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3694 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3693 47 43 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3692 43 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3691 12 12 43 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3690 43 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M3689 43 44 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D3687 are shorted:
* D3687 12 12 D_lateral AREA=3.75E-016    ; (-1695.501 200 -1695.5 206)CMOSN3687 12 12 D_lateral AREA=3.75E-016    
* Pins of element D3686 are shorted:
* D3686 12 12 D_lateral AREA=2f    ; (-1714.5 197 -1704.499 209)CMOSN3686 12 12 D_lateral AREA=2f    
* Pins of element D3685 are shorted:
* D3685 12 12 D_lateral AREA=2.3749375f    ; (-1760.5 232 -1726.5 236)CMOSN3685 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3684 are shorted:
* D3684 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 248 -1760.499 252)CMOSN3684 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3683 are shorted:
* D3683 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 264 -1760.499 268)CMOSN3683 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3682 are shorted:
* D3682 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 280 -1760.499 284)CMOSN3682 12 12 D_lateral AREA=2.5E-016    
M3674 8 46 45 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3673 45 46 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3672 8 46 45 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3671 45 46 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3670 8 46 45 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3669 45 46 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3668 46 47 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3667 46 47 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M3666 44 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D3664 are shorted:
* D3664 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 110 -1605.499 114)CMOSN3664 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3663 are shorted:
* D3663 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 126 -1605.499 130)CMOSN3663 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3662 are shorted:
* D3662 8 8 D_lateral AREA=8.625f    ; (-1668.5 142 -1605.499 154)CMOSN3662 8 8 D_lateral AREA=8.625f    
* Pins of element D3661 are shorted:
* D3661 8 8 D_lateral AREA=4.375E-016    ; (-1673.501 146 -1673.5 153)CMOSN3661 8 8 D_lateral AREA=4.375E-016    
* Pins of element D3660 are shorted:
* D3660 8 8 D_lateral AREA=4.1250625f    ; (-1673.501 166 -1615.5 174.001)CMOSN3660 8 8 D_lateral AREA=4.1250625f    
* Pins of element D3659 are shorted:
* D3659 8 8 D_lateral AREA=4.062625f    ; (-1674.501 183.999 -1621.499 190)CMOSN3659 8 8 D_lateral AREA=4.062625f    
M3658 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3657 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3656 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3655 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3654 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3653 45 46 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3652 44 12 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M3651 46 47 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M3650 46 47 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D3649 are shorted:
* D3649 12 12 D_lateral AREA=2.4374375f    ; (-1730.5 166 -1697.5 172)CMOSN3649 12 12 D_lateral AREA=2.4374375f    
* Pins of element D3648 are shorted:
* D3648 12 12 D_lateral AREA=2.687375f    ; (-1732.5 150 -1697.5 154)CMOSN3648 12 12 D_lateral AREA=2.687375f    
* Pins of element D3646 are shorted:
* D3646 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 110 -1733.499 114)CMOSN3646 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3645 are shorted:
* D3645 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 126 -1733.499 130)CMOSN3645 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3644 are shorted:
* D3644 12 12 D_lateral AREA=2.3749375f    ; (-1733.5 142 -1699.5 146)CMOSN3644 12 12 D_lateral AREA=2.3749375f    
C3637 12 12  184.041f    ; (1836.5 85 2122.5 371)CMOSN.041f    
M3636 45 46 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
* Pins of element D3635 are shorted:
* D3635 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 94 -1605.499 98)CMOSN3635 8 8 D_lateral AREA=2.5E-016    
M3634 45 46 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
* Pins of element D3633 are shorted:
* D3633 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 94 -1733.499 98)CMOSN3633 12 12 D_lateral AREA=2.5E-016    
C3630 47 12  184.041f    ; (-2185.5 85 -1899.5 371)CMOSN.041f    
M3620 48 52 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3619 48 52 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3618 48 52 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D3617 are shorted:
* D3617 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -96 1697.5 -92)CMOSN3617 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3616 are shorted:
* D3616 12 12 D_lateral AREA=3.249875f    ; (1661.5 -80 1697.5 -72)CMOSN3616 12 12 D_lateral AREA=3.249875f    
* Pins of element D3614 are shorted:
* D3614 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -93 1637.501 -89)CMOSN3614 8 8 D_lateral AREA=2.5E-016    
M3612 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3610 48 50 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3608 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3606 48 50 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3603 48 50 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3602 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3601 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3600 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D3599 are shorted:
* D3599 8 8 D_lateral AREA=8.875125f    ; (1502.499 -77 1637.501 -72.999)CMOSN3599 8 8 D_lateral AREA=8.875125f    
M3593 8 49 59 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3591 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3589 8 49 59 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3587 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3584 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3583 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3582 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3581 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3580 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3579 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3578 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3577 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D3575 are shorted:
* D3575 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -92 -1760.499 -88)CMOSN3575 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3574 are shorted:
* D3574 12 12 D_lateral AREA=3.249875f    ; (-1760.5 -76 -1724.5 -68)CMOSN3574 12 12 D_lateral AREA=3.249875f    
* Pins of element D3573 are shorted:
* D3573 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -105 -1700.5 -101)CMOSN3573 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3572 are shorted:
* D3572 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -89 -1700.5 -85)CMOSN3572 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3571 are shorted:
* D3571 8 8 D_lateral AREA=8.875125f    ; (-1700.501 -73 -1565.499 -68.999)CMOSN3571 8 8 D_lateral AREA=8.875125f    
M3559 50 8 52 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M3558 52 8 50 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M3557 50 8 52 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M3556 12 52 48 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M3555 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3554 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3553 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3552 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3551 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3550 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3549 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3548 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3547 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3546 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3545 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3544 12 52 48 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
* Pins of element D3541 are shorted:
* D3541 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -192 1697.5 -188)CMOSN3541 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3540 are shorted:
* D3540 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -176 1697.5 -172)CMOSN3540 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3539 are shorted:
* D3539 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -160 1697.5 -156)CMOSN3539 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3538 are shorted:
* D3538 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -144 1697.5 -140)CMOSN3538 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3537 are shorted:
* D3537 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -128 1697.5 -124)CMOSN3537 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3536 are shorted:
* D3536 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -112 1697.5 -108)CMOSN3536 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3535 are shorted:
* D3535 8 8 D_lateral AREA=1.8125625f    ; (1614.5 -143.001 1637.501 -137)CMOSN3535 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3534 are shorted:
* D3534 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -125 1637.501 -121)CMOSN3534 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3533 are shorted:
* D3533 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -109 1637.501 -105)CMOSN3533 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3532 are shorted:
* D3532 8 8 D_lateral AREA=3.125E-016    ; (1611.5 -201 1611.501 -196)CMOSN3532 8 8 D_lateral AREA=3.125E-016    
M3531 50 72 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M3530 50 72 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M3529 50 72 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M3528 50 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M3527 8 50 48 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3525 48 50 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3523 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3521 48 50 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D3519 are shorted:
* D3519 8 8 D_lateral AREA=3.125E-016    ; (1558.499 -201 1558.5 -196)CMOSN3519 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3518 are shorted:
* D3518 8 8 D_lateral AREA=2.5E-016    ; (1558.499 -184 1558.5 -180)CMOSN3518 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3517 are shorted:
* D3517 8 8 D_lateral AREA=3.5625625f    ; (1558.499 -168 1605.5 -157.999)CMOSN3517 8 8 D_lateral AREA=3.5625625f    
M3516 8 50 48 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3515 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3514 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3513 8 50 48 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3508 8 12 49 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M3507 49 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M3506 49 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M3505 49 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M3504 8 49 59 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3502 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3500 8 49 59 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3498 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
* Pins of element D3495 are shorted:
* D3495 8 8 D_lateral AREA=2.5E-016    ; (-1621.5 -180 -1621.499 -176)CMOSN3495 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3494 are shorted:
* D3494 8 8 D_lateral AREA=3.5625625f    ; (-1668.5 -164 -1621.499 -153.999)CMOSN3494 8 8 D_lateral AREA=3.5625625f    
* Pins of element D3493 are shorted:
* D3493 8 8 D_lateral AREA=3.125E-016    ; (-1621.5 -197 -1621.499 -192)CMOSN3493 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3492 are shorted:
* D3492 8 8 D_lateral AREA=3.125E-016    ; (-1674.501 -197 -1674.5 -192)CMOSN3492 8 8 D_lateral AREA=3.125E-016    
M3491 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M3490 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3489 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3488 59 49 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3487 56 12 49 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M3486 49 12 56 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M3485 56 12 49 12 CMOSN L=500n W=3.25u AD=2.53125p PD=5u AS=4.875p PS=9.5u    
M3484 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3483 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3482 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3481 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3480 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3479 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3478 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3477 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3476 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3475 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3474 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3473 59 56 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3472 56 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
* Pins of element D3471 are shorted:
* D3471 12 12 D_lateral AREA=2.3749375f    ; (-1760.5 -204 -1726.5 -200)CMOSN3471 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3470 are shorted:
* D3470 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -188 -1760.499 -184)CMOSN3470 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3469 are shorted:
* D3469 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -172 -1760.499 -168)CMOSN3469 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3468 are shorted:
* D3468 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -156 -1760.499 -152)CMOSN3468 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3467 are shorted:
* D3467 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -140 -1760.499 -136)CMOSN3467 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3466 are shorted:
* D3466 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -124 -1760.499 -120)CMOSN3466 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3465 are shorted:
* D3465 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -108 -1760.499 -104)CMOSN3465 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3464 are shorted:
* D3464 8 8 D_lateral AREA=1.8125625f    ; (-1700.501 -139.001 -1677.5 -133)CMOSN3464 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3463 are shorted:
* D3463 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -121 -1700.5 -117)CMOSN3463 8 8 D_lateral AREA=2.5E-016    
M3455 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3454 52 72 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3453 12 72 52 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3452 52 72 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M3451 52 53 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M3450 53 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M3449 51 48 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M3448 51 48 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D3447 are shorted:
* D3447 12 12 D_lateral AREA=2f    ; (1641.499 -243 1651.5 -231)CMOSN3447 12 12 D_lateral AREA=2f    
* Pins of element D3446 are shorted:
* D3446 12 12 D_lateral AREA=2.687375f    ; (1634.5 -290 1669.5 -286)CMOSN3446 12 12 D_lateral AREA=2.687375f    
* Pins of element D3445 are shorted:
* D3445 12 12 D_lateral AREA=2.4374375f    ; (1634.5 -274 1667.5 -268)CMOSN3445 12 12 D_lateral AREA=2.4374375f    
* Pins of element D3444 are shorted:
* D3444 12 12 D_lateral AREA=2.3749375f    ; (1663.5 -208 1697.5 -204)CMOSN3444 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3443 are shorted:
* D3443 12 12 D_lateral AREA=2.3749375f    ; (1636.5 -298 1670.5 -294)CMOSN3443 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3442 are shorted:
* D3442 12 12 D_lateral AREA=3.75E-016    ; (1632.5 -240 1632.501 -234)CMOSN3442 12 12 D_lateral AREA=3.75E-016    
M3440 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3439 51 48 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3438 51 48 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M3437 52 53 50 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M3436 50 53 52 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3435 52 53 50 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M3434 53 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D3433 are shorted:
* D3433 8 8 D_lateral AREA=4.1250625f    ; (1552.5 -274 1610.501 -265.999)CMOSN3433 8 8 D_lateral AREA=4.1250625f    
* Pins of element D3432 are shorted:
* D3432 8 8 D_lateral AREA=4.375E-016    ; (1610.5 -294 1610.501 -287)CMOSN3432 8 8 D_lateral AREA=4.375E-016    
* Pins of element D3431 are shorted:
* D3431 8 8 D_lateral AREA=8.625f    ; (1542.499 -298 1605.5 -286)CMOSN3431 8 8 D_lateral AREA=8.625f    
* Pins of element D3430 are shorted:
* D3430 8 8 D_lateral AREA=4.062625f    ; (1558.499 -256.001 1611.501 -250)CMOSN3430 8 8 D_lateral AREA=4.062625f    
M3429 8 58 54 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3428 54 58 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3427 58 59 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M3426 58 59 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M3425 56 55 49 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M3424 49 55 56 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3423 56 55 49 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M3422 55 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D3421 are shorted:
* D3421 8 8 D_lateral AREA=8.625f    ; (-1668.5 -294 -1605.499 -282)CMOSN3421 8 8 D_lateral AREA=8.625f    
* Pins of element D3420 are shorted:
* D3420 8 8 D_lateral AREA=4.375E-016    ; (-1673.501 -290 -1673.5 -283)CMOSN3420 8 8 D_lateral AREA=4.375E-016    
* Pins of element D3419 are shorted:
* D3419 8 8 D_lateral AREA=4.1250625f    ; (-1673.501 -270 -1615.5 -261.999)CMOSN3419 8 8 D_lateral AREA=4.1250625f    
* Pins of element D3418 are shorted:
* D3418 8 8 D_lateral AREA=4.062625f    ; (-1674.501 -252.001 -1621.499 -246)CMOSN3418 8 8 D_lateral AREA=4.062625f    
M3417 12 58 54 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3416 54 58 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3415 56 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3414 12 12 56 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3413 56 55 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M3412 55 12 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M3411 58 59 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M3410 58 59 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D3409 are shorted:
* D3409 12 12 D_lateral AREA=3.75E-016    ; (-1695.501 -236 -1695.5 -230)CMOSN3409 12 12 D_lateral AREA=3.75E-016    
* Pins of element D3408 are shorted:
* D3408 12 12 D_lateral AREA=2f    ; (-1714.5 -239 -1704.499 -227)CMOSN3408 12 12 D_lateral AREA=2f    
* Pins of element D3407 are shorted:
* D3407 12 12 D_lateral AREA=2.4374375f    ; (-1730.5 -270 -1697.5 -264)CMOSN3407 12 12 D_lateral AREA=2.4374375f    
* Pins of element D3406 are shorted:
* D3406 12 12 D_lateral AREA=2.687375f    ; (-1732.5 -286 -1697.5 -282)CMOSN3406 12 12 D_lateral AREA=2.687375f    
* Pins of element D3405 are shorted:
* D3405 12 12 D_lateral AREA=2.3749375f    ; (-1733.5 -294 -1699.5 -290)CMOSN3405 12 12 D_lateral AREA=2.3749375f    
C3398 48 12  184.041f    ; (1836.5 -355 2122.5 -69)CMOSN.041f    
M3397 57 51 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M3396 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3395 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3394 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3393 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3392 57 51 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D3391 are shorted:
* D3391 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -346 1670.5 -342)CMOSN3391 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3390 are shorted:
* D3390 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -330 1670.5 -326)CMOSN3390 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3389 are shorted:
* D3389 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -314 1670.5 -310)CMOSN3389 12 12 D_lateral AREA=2.5E-016    
M3388 57 51 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M3387 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3386 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3385 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3384 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3383 57 51 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
* Pins of element D3382 are shorted:
* D3382 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -346 1542.5 -342)CMOSN3382 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3381 are shorted:
* D3381 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -330 1542.5 -326)CMOSN3381 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3380 are shorted:
* D3380 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -314 1542.5 -310)CMOSN3380 8 8 D_lateral AREA=2.5E-016    
M3379 54 58 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M3378 8 58 54 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3377 54 58 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M3376 8 58 54 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M3375 54 58 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
* Pins of element D3374 are shorted:
* D3374 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -342 -1605.499 -338)CMOSN3374 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3373 are shorted:
* D3373 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -326 -1605.499 -322)CMOSN3373 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3372 are shorted:
* D3372 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -310 -1605.499 -306)CMOSN3372 8 8 D_lateral AREA=2.5E-016    
M3371 54 58 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M3370 54 58 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3369 54 58 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3368 54 58 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3367 54 58 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D3366 are shorted:
* D3366 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -342 -1733.499 -338)CMOSN3366 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3365 are shorted:
* D3365 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -326 -1733.499 -322)CMOSN3365 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3364 are shorted:
* D3364 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -310 -1733.499 -306)CMOSN3364 12 12 D_lateral AREA=2.5E-016    
C3361 59 12  184.041f    ; (-2185.5 -351 -1899.5 -65)CMOSN.041f    
M3336 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3335 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3334 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3333 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3332 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3331 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3330 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3329 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3328 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3327 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3326 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D3325 are shorted:
* D3325 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -596 1697.5 -592)CMOSN3325 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3324 are shorted:
* D3324 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -580 1697.5 -576)CMOSN3324 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3323 are shorted:
* D3323 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -564 1697.5 -560)CMOSN3323 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3322 are shorted:
* D3322 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -548 1697.5 -544)CMOSN3322 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3321 are shorted:
* D3321 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -532 1697.5 -528)CMOSN3321 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3320 are shorted:
* D3320 12 12 D_lateral AREA=3.249875f    ; (1661.5 -516 1697.5 -508)CMOSN3320 12 12 D_lateral AREA=3.249875f    
* Pins of element D3319 are shorted:
* D3319 8 8 D_lateral AREA=1.8125625f    ; (1614.5 -579.001 1637.501 -573)CMOSN3319 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3318 are shorted:
* D3318 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -561 1637.501 -557)CMOSN3318 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3317 are shorted:
* D3317 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -545 1637.501 -541)CMOSN3317 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3316 are shorted:
* D3316 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -529 1637.501 -525)CMOSN3316 8 8 D_lateral AREA=2.5E-016    
M3313 8 61 60 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3311 60 61 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3309 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3307 60 61 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3305 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3303 60 61 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3301 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3299 60 61 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
* Pins of element D3296 are shorted:
* D3296 8 8 D_lateral AREA=3.5625625f    ; (1558.499 -604 1605.5 -593.999)CMOSN3296 8 8 D_lateral AREA=3.5625625f    
M3295 60 61 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3294 8 61 60 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3293 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3292 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3291 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3290 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3289 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3288 8 61 60 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D3287 are shorted:
* D3287 8 8 D_lateral AREA=8.875125f    ; (1502.499 -513 1637.501 -508.999)CMOSN3287 8 8 D_lateral AREA=8.875125f    
M3285 8 73 70 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3284 70 45 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3283 are shorted:
* D3283 8 8 D_lateral AREA=3.125E-016    ; (701.5 -603.5 701.501 -598.5)CMOSN3283 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3281 are shorted:
* D3281 8 8 D_lateral AREA=3.125E-016    ; (417 -603.5 417.001 -598.5)CMOSN3281 8 8 D_lateral AREA=3.125E-016    
M3280 8 83 84 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3279 84 45 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3277 8 18 91 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3276 91 45 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3275 are shorted:
* D3275 8 8 D_lateral AREA=3.125E-016    ; (133 -603.5 133.001 -598.5)CMOSN3275 8 8 D_lateral AREA=3.125E-016    
M3273 8 334 101 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3272 101 45 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3271 are shorted:
* D3271 8 8 D_lateral AREA=3.125E-016    ; (-151.5 -603.5 -151.499 -598.5)CMOSN3271 8 8 D_lateral AREA=3.125E-016    
M3258 8 40 128 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3257 128 45 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
* Pins of element D3256 are shorted:
* D3256 8 8 D_lateral AREA=3.125E-016    ; (-733 -604.5 -732.999 -599.5)CMOSN3256 8 8 D_lateral AREA=3.125E-016    
M3236 150 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M3235 8 150 249 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M3233 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3231 8 150 249 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3229 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3227 8 150 249 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3225 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3223 8 150 249 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M3221 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
* Pins of element D3218 are shorted:
* D3218 8 8 D_lateral AREA=3.5625625f    ; (-1668.5 -600 -1621.499 -589.999)CMOSN3218 8 8 D_lateral AREA=3.5625625f    
M3217 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M3216 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3215 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3214 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3213 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3212 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3211 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M3210 249 150 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M3209 148 12 150 12 CMOSN L=500n W=3.25u AD=2.53125p PD=5u AS=4.875p PS=9.5u    
M3208 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3207 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3206 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3205 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3204 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3203 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3202 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3201 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3200 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3199 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3198 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3197 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D3196 are shorted:
* D3196 12 12 D_lateral AREA=3.249875f    ; (-1760.5 -512 -1724.5 -504)CMOSN3196 12 12 D_lateral AREA=3.249875f    
* Pins of element D3194 are shorted:
* D3194 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -592 -1760.499 -588)CMOSN3194 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3193 are shorted:
* D3193 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -576 -1760.499 -572)CMOSN3193 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3192 are shorted:
* D3192 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -560 -1760.499 -556)CMOSN3192 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3191 are shorted:
* D3191 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -544 -1760.499 -540)CMOSN3191 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3190 are shorted:
* D3190 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -528 -1760.499 -524)CMOSN3190 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3188 are shorted:
* D3188 8 8 D_lateral AREA=1.8125625f    ; (-1700.501 -575.001 -1677.5 -569)CMOSN3188 8 8 D_lateral AREA=1.8125625f    
* Pins of element D3187 are shorted:
* D3187 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -557 -1700.5 -553)CMOSN3187 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3186 are shorted:
* D3186 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -541 -1700.5 -537)CMOSN3186 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3185 are shorted:
* D3185 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -525 -1700.5 -521)CMOSN3185 8 8 D_lateral AREA=2.5E-016    
* Pins of element D3184 are shorted:
* D3184 8 8 D_lateral AREA=8.875125f    ; (-1700.501 -509 -1565.499 -504.999)CMOSN3184 8 8 D_lateral AREA=8.875125f    
M3176 61 8 63 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M3175 63 8 61 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M3174 61 8 63 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M3173 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M3172 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3171 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3170 60 63 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M3169 12 63 60 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M3168 63 160 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3167 12 160 63 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M3166 63 160 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M3165 63 64 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M3164 64 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
* Pins of element D3163 are shorted:
* D3163 12 12 D_lateral AREA=2f    ; (1641.499 -679 1651.5 -667)CMOSN3163 12 12 D_lateral AREA=2f    
* Pins of element D3161 are shorted:
* D3161 12 12 D_lateral AREA=2.3749375f    ; (1663.5 -644 1697.5 -640)CMOSN3161 12 12 D_lateral AREA=2.3749375f    
* Pins of element D3160 are shorted:
* D3160 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -628 1697.5 -624)CMOSN3160 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3159 are shorted:
* D3159 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -612 1697.5 -608)CMOSN3159 12 12 D_lateral AREA=2.5E-016    
* Pins of element D3158 are shorted:
* D3158 12 12 D_lateral AREA=3.75E-016    ; (1632.5 -676 1632.501 -670)CMOSN3158 12 12 D_lateral AREA=3.75E-016    
* Pins of element D3156 are shorted:
* D3156 8 8 D_lateral AREA=3.125E-016    ; (1611.5 -637 1611.501 -632)CMOSN3156 8 8 D_lateral AREA=3.125E-016    
M3155 61 160 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M3154 61 160 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M3153 61 160 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M3152 63 64 61 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M3151 61 64 63 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M3150 63 64 61 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M3149 64 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M3148 61 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
* Pins of element D3146 are shorted:
* D3146 8 8 D_lateral AREA=4.062625f    ; (1558.499 -692.001 1611.501 -686)CMOSN3146 8 8 D_lateral AREA=4.062625f    
* Pins of element D3145 are shorted:
* D3145 8 8 D_lateral AREA=3.125E-016    ; (1558.499 -637 1558.5 -632)CMOSN3145 8 8 D_lateral AREA=3.125E-016    
* Pins of element D3144 are shorted:
* D3144 8 8 D_lateral AREA=2.5E-016    ; (1558.499 -620 1558.5 -616)CMOSN3144 8 8 D_lateral AREA=2.5E-016    
M3143 8 69 66 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3142 66 65 163 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3141 65 82 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3140 8 82 68 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3139 68 69 160 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M3138 68 65 160 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3137 12 69 163 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3136 163 65 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3135 65 82 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M3134 67 82 160 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M3133 160 69 67 12 CMOSN L=750n W=750n AD=7.375p PD=19u AS=968.75f PS=3u    
M3132 12 65 67 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M3131 8 70 72 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3130 68 161 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3129 8 161 69 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3128 161 71 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3127 12 70 72 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3126 67 161 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3125 12 161 69 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3124 161 71 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3120 8 73 71 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M3119 71 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M3118 70 73 75 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3117 75 45 12 12 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3116 74 54 71 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M3115 12 73 74 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D3114 are shorted:
* D3114 12 12 D_lateral AREA=3.125E-016    ; (709 -702 714 -701.999)CMOSN3114 12 12 D_lateral AREA=3.125E-016    
M3113 8 80 79 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3112 79 76 175 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3111 76 94 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3110 8 94 78 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3109 78 80 172 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M3108 78 173 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3107 78 76 172 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3106 12 80 175 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3105 175 76 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3104 76 94 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M3103 77 94 172 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M3102 77 80 172 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M3101 77 173 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3100 12 76 77 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M3099 8 84 82 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3098 8 173 80 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3097 173 85 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3096 12 84 82 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3095 12 173 80 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3094 173 85 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3093 81 54 85 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M3092 12 83 81 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D3091 are shorted:
* D3091 12 12 D_lateral AREA=3.125E-016    ; (424.5 -702 429.5 -701.999)CMOSN3091 12 12 D_lateral AREA=3.125E-016    
M3090 8 83 85 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M3089 85 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M3088 8 180 87 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3087 87 88 182 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3086 84 83 86 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3085 86 45 12 12 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3084 12 180 182 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3083 182 88 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3082 88 104 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3081 8 104 90 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3080 90 189 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3079 8 189 180 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3078 90 180 188 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M3077 90 88 188 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3076 88 104 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M3075 89 104 188 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M3074 89 189 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3073 12 189 180 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3072 89 180 188 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M3071 12 88 89 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M3070 8 91 94 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3069 189 95 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3068 12 91 94 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3067 91 18 93 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3066 93 45 12 12 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3065 189 95 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3064 92 54 95 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M3063 12 18 92 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D3062 are shorted:
* D3062 12 12 D_lateral AREA=3.125E-016    ; (140.5 -702 145.5 -701.999)CMOSN3062 12 12 D_lateral AREA=3.125E-016    
M3061 8 18 95 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M3060 95 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M3059 8 100 96 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3058 96 99 197 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3057 12 100 197 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3056 197 99 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3055 99 116 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3054 8 116 98 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3053 98 202 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3052 8 202 100 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3051 98 100 192 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M3050 98 99 192 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3049 99 116 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M3048 97 116 192 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M3047 97 202 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3046 12 202 100 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3045 97 100 192 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M3044 12 99 97 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M3043 8 101 104 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M3042 202 105 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M3041 8 334 105 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M3040 12 101 104 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M3039 101 334 103 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3038 103 45 12 12 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3037 202 105 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M3036 102 54 105 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M3035 12 334 102 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D3034 are shorted:
* D3034 12 12 D_lateral AREA=3.125E-016    ; (-144 -702 -139 -701.999)CMOSN3034 12 12 D_lateral AREA=3.125E-016    
M3033 8 117 109 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3032 109 118 108 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M3031 105 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M3029 107 114 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M3028 203 215 107 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M3027 8 119 106 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3025 12 117 108 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3024 108 118 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3023 203 114 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M3022 12 215 203 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M3021 12 119 114 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M3020 118 8 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3019 8 62 115 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M3018 8 62 117 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3017 116 117 115 8 CMOSP L=750n W=750n AD=7.4375p PD=19.125u AS=968.75f PS=3u    
M3016 115 118 116 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3015 8 8 115 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3014 114 111 106 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M3013 111 108 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M3012 8 108 113 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M3011 113 119 222 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M3010 113 120 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3009 8 120 119 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3008 113 111 222 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M3007 118 8 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M3006 110 8 116 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M3005 110 62 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M3004 12 62 117 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M3003 110 117 116 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M3002 12 118 110 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M3001 114 111 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M3000 111 108 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2999 112 108 222 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2998 112 119 222 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2997 112 120 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2996 12 120 119 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2995 12 111 112 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2994 62 121 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2993 8 37 121 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2992 8 221 120 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2990 62 121 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2989 122 45 121 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2988 12 37 122 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2987 12 221 120 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
* Pins of element D2986 are shorted:
* D2986 12 12 D_lateral AREA=3.125E-016    ; (-441 -624 -436 -623.999)CMOSN2986 12 12 D_lateral AREA=3.125E-016    
M2985 121 45 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2984 8 127 123 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2983 123 126 232 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2982 8 143 126 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2980 12 127 232 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2979 232 126 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2978 12 143 126 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2977 125 130 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2976 8 130 127 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2975 125 127 228 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2974 125 126 228 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2973 8 143 125 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2972 124 130 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2971 12 130 127 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2970 124 127 228 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2969 12 126 124 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2968 124 143 228 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2967 8 128 132 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2966 130 235 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M2965 8 40 235 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2964 235 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2963 12 128 132 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2962 128 40 131 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2961 131 45 12 12 CMOSN L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2960 130 235 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M2959 129 54 235 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2958 12 40 129 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2957 are shorted:
* D2957 12 12 D_lateral AREA=3.125E-016    ; (-725.5 -703 -720.5 -702.999)CMOSN2957 12 12 D_lateral AREA=3.125E-016    
M2956 8 141 134 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2955 134 137 244 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2954 8 142 133 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2953 133 140 242 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2952 12 141 244 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2951 244 137 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2950 12 142 242 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2949 242 140 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2948 137 242 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2947 8 242 136 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2946 136 144 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2945 8 144 141 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2944 136 141 238 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2943 136 137 238 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2942 140 8 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2941 8 146 139 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2940 8 146 142 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2939 143 142 139 8 CMOSP L=750n W=750n AD=7.4375p PD=19.125u AS=968.75f PS=3u    
M2938 139 140 143 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2937 8 8 139 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2936 137 242 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2935 135 242 238 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2934 135 144 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2933 12 144 141 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2932 135 141 238 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2931 12 137 135 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2930 140 8 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2929 138 8 143 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2928 138 146 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2927 12 146 142 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2926 138 142 143 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2925 12 140 138 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2924 8 41 144 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2923 144 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2922 8 41 146 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2921 146 45 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2920 147 54 144 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2919 12 41 147 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2918 145 45 146 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2917 12 41 145 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2916 are shorted:
* D2916 12 12 D_lateral AREA=3.125E-016    ; (-1002.5 -703 -997.5 -702.999)CMOSN2916 12 12 D_lateral AREA=3.125E-016    
* Pins of element D2915 are shorted:
* D2915 12 12 D_lateral AREA=3.125E-016    ; (-1002.5 -625 -997.5 -624.999)CMOSN2915 12 12 D_lateral AREA=3.125E-016    
M2914 8 12 150 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M2913 150 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M2912 150 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M2911 148 149 150 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M2910 150 149 148 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M2909 148 149 150 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M2908 149 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D2906 are shorted:
* D2906 8 8 D_lateral AREA=4.062625f    ; (-1674.501 -688.001 -1621.499 -682)CMOSN2906 8 8 D_lateral AREA=4.062625f    
* Pins of element D2905 are shorted:
* D2905 8 8 D_lateral AREA=2.5E-016    ; (-1621.5 -616 -1621.499 -612)CMOSN2905 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2904 are shorted:
* D2904 8 8 D_lateral AREA=3.125E-016    ; (-1621.5 -633 -1621.499 -628)CMOSN2904 8 8 D_lateral AREA=3.125E-016    
* Pins of element D2903 are shorted:
* D2903 8 8 D_lateral AREA=3.125E-016    ; (-1674.501 -633 -1674.5 -628)CMOSN2903 8 8 D_lateral AREA=3.125E-016    
M2902 148 12 150 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M2901 150 12 148 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M2900 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M2899 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2898 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2897 249 148 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2896 148 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M2895 12 12 148 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M2894 148 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M2893 148 149 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M2892 149 12 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
* Pins of element D2891 are shorted:
* D2891 12 12 D_lateral AREA=3.75E-016    ; (-1695.501 -672 -1695.5 -666)CMOSN2891 12 12 D_lateral AREA=3.75E-016    
* Pins of element D2890 are shorted:
* D2890 12 12 D_lateral AREA=2f    ; (-1714.5 -675 -1704.499 -663)CMOSN2890 12 12 D_lateral AREA=2f    
* Pins of element D2888 are shorted:
* D2888 12 12 D_lateral AREA=2.3749375f    ; (-1760.5 -640 -1726.5 -636)CMOSN2888 12 12 D_lateral AREA=2.3749375f    
* Pins of element D2887 are shorted:
* D2887 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -624 -1760.499 -620)CMOSN2887 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2886 are shorted:
* D2886 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -608 -1760.499 -604)CMOSN2886 12 12 D_lateral AREA=2.5E-016    
C2879 60 12  184.041f    ; (1836.5 -791 2122.5 -505)CMOSN.041f    
M2878 152 151 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M2877 12 151 152 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M2876 152 151 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2875 12 151 152 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M2874 152 151 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2873 12 151 152 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M2872 152 151 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M2871 151 60 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M2870 151 60 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D2869 are shorted:
* D2869 12 12 D_lateral AREA=2.687375f    ; (1634.5 -726 1669.5 -722)CMOSN2869 12 12 D_lateral AREA=2.687375f    
* Pins of element D2868 are shorted:
* D2868 12 12 D_lateral AREA=2.4374375f    ; (1634.5 -710 1667.5 -704)CMOSN2868 12 12 D_lateral AREA=2.4374375f    
* Pins of element D2867 are shorted:
* D2867 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -782 1670.5 -778)CMOSN2867 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2866 are shorted:
* D2866 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -766 1670.5 -762)CMOSN2866 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2865 are shorted:
* D2865 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -750 1670.5 -746)CMOSN2865 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2864 are shorted:
* D2864 12 12 D_lateral AREA=2.3749375f    ; (1636.5 -734 1670.5 -730)CMOSN2864 12 12 D_lateral AREA=2.3749375f    
M2863 152 151 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M2862 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2861 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2860 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2859 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2858 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2857 152 151 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M2856 151 60 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M2855 151 60 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
* Pins of element D2854 are shorted:
* D2854 8 8 D_lateral AREA=4.1250625f    ; (1552.5 -710 1610.501 -701.999)CMOSN2854 8 8 D_lateral AREA=4.1250625f    
* Pins of element D2853 are shorted:
* D2853 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -782 1542.5 -778)CMOSN2853 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2852 are shorted:
* D2852 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -766 1542.5 -762)CMOSN2852 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2851 are shorted:
* D2851 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -750 1542.5 -746)CMOSN2851 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2850 are shorted:
* D2850 8 8 D_lateral AREA=4.375E-016    ; (1610.5 -730 1610.501 -723)CMOSN2850 8 8 D_lateral AREA=4.375E-016    
* Pins of element D2849 are shorted:
* D2849 8 8 D_lateral AREA=8.625f    ; (1542.499 -734 1605.5 -722)CMOSN2849 8 8 D_lateral AREA=8.625f    
M2848 8 251 267 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2847 156 153 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2846 251 252 156 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2845 155 253 252 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2844 8 264 155 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2842 8 162 154 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2841 154 159 153 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2839 251 153 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2838 12 252 251 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2837 12 162 153 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2836 153 159 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2834 8 263 264 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2833 8 172 253 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2832 8 172 266 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2831 266 253 265 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2830 266 264 265 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2829 266 263 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2828 8 163 159 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2827 8 163 158 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2826 158 164 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2825 8 164 162 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2824 158 162 263 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2823 158 159 263 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2822 12 163 159 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2821 157 163 263 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2820 157 164 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2819 12 164 162 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2818 157 162 263 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2817 12 159 157 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2816 8 165 164 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2813 272 274 166 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2811 12 165 164 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2809 12 274 272 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2807 8 272 288 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2806 8 167 166 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=562.5f PS=2.25u    
M2805 169 275 274 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2804 8 284 169 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2803 8 188 275 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2802 8 188 286 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2801 8 174 168 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2800 168 176 167 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2799 176 175 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2798 8 175 171 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2797 12 167 272 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=968.75f PS=3u    
M2796 12 174 167 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2795 167 176 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2794 176 175 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2793 12 176 170 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2792 8 290 177 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2791 8 283 284 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2790 286 275 285 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2789 286 284 285 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2788 286 283 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2787 171 177 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2786 8 177 174 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2785 171 174 283 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2784 171 176 283 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2783 12 290 177 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2781 170 177 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2780 12 177 174 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2779 170 174 283 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2778 170 175 283 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2775 8 291 295 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2774 178 181 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2773 291 297 178 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2772 291 181 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2771 12 297 291 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2770 184 298 297 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2769 8 309 184 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2768 8 192 298 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2767 8 192 311 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2766 311 298 310 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2765 8 190 183 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2764 183 179 181 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2763 179 182 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2762 8 182 186 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2761 186 179 308 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2760 12 190 181 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2759 181 179 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2758 179 182 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2757 185 182 308 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2756 12 179 185 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2755 8 307 187 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2754 8 308 309 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2753 311 309 310 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2752 311 308 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2751 186 187 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2750 8 187 190 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2749 186 190 308 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2748 12 307 187 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2746 185 187 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2745 12 187 190 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2744 185 190 308 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2741 8 313 320 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2740 191 196 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2739 313 322 191 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2738 313 196 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2737 12 322 313 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2736 199 324 322 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2735 8 332 199 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2734 8 220 324 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2733 8 220 323 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2732 323 324 329 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2731 323 332 329 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2729 8 200 198 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2728 198 193 196 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2727 193 197 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2726 8 197 195 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2725 195 200 331 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2723 195 193 331 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2722 12 200 196 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2721 196 193 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2720 193 197 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2719 194 197 331 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2718 194 200 331 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2716 12 193 194 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2715 8 330 201 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2714 8 331 332 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2713 8 331 323 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2712 8 201 195 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2711 8 201 200 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2710 12 330 201 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2708 12 201 194 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2707 12 201 200 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2706 8 203 214 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2705 8 217 207 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2701 8 335 344 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2700 206 216 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2699 335 346 206 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2697 8 350 205 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2696 8 218 204 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2694 12 203 214 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2693 12 217 215 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2692 335 216 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2691 12 346 335 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2690 12 218 216 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2689 215 208 207 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2688 208 132 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2687 220 217 210 8 CMOSP L=750n W=750n AD=7.4375p PD=19.125u AS=968.75f PS=3u    
M2686 8 222 210 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2685 8 222 217 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2684 210 208 220 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2683 8 132 210 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2682 346 348 205 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2681 8 353 350 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2680 8 228 348 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2679 8 228 347 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2678 347 348 354 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2677 347 350 354 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2676 347 353 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2675 216 211 204 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2674 211 214 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2673 8 214 213 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2672 213 218 353 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2671 213 219 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2670 8 219 218 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2669 213 211 353 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2668 215 208 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2667 208 132 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2666 209 132 220 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2665 209 217 220 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2664 209 222 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2663 12 222 217 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2662 12 208 209 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2661 216 211 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2660 211 214 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2659 212 214 353 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2658 212 218 353 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2657 212 219 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2656 12 219 218 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2655 12 211 212 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2654 8 37 221 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2653 8 352 219 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2651 223 54 221 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2650 12 37 223 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2649 12 352 219 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
* Pins of element D2647 are shorted:
* D2647 12 12 D_lateral AREA=3.125E-016    ; (-441 -727 -436 -726.999)CMOSN2647 12 12 D_lateral AREA=3.125E-016    
M2646 221 54 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2644 8 357 367 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2643 227 224 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2642 357 358 227 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2641 226 371 358 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2640 8 369 226 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2639 8 233 225 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2638 225 229 224 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2637 357 224 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2636 12 358 357 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2635 12 233 224 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2634 224 229 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2633 8 236 369 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2632 8 238 371 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2631 8 238 370 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2630 370 371 373 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2629 370 369 373 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2628 370 236 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2627 229 232 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2626 8 232 231 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2625 231 234 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2624 8 234 233 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2623 231 233 236 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2622 231 229 236 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2621 229 232 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2620 230 232 236 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2619 230 234 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2618 12 234 233 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2617 230 233 236 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2616 12 229 230 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2615 8 375 234 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2612 12 375 234 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2610 8 243 237 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2609 237 241 383 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2608 12 243 383 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2607 383 241 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2606 241 244 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2605 8 244 240 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2604 240 245 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2603 8 245 243 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2602 240 243 381 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2601 240 241 381 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2600 241 244 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2599 239 244 381 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2598 239 245 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2597 12 245 243 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2596 239 243 381 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2595 12 241 239 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2594 8 41 245 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2593 245 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2592 246 248 245 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2591 12 41 246 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2590 are shorted:
* D2590 12 12 D_lateral AREA=3.125E-016    ; (-1002.5 -798 -997.5 -797.999)CMOSN2590 12 12 D_lateral AREA=3.125E-016    
M2589 248 247 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M2588 8 247 248 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M2587 248 247 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2586 8 247 248 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M2585 248 247 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M2584 8 247 248 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M2583 248 247 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M2582 247 249 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M2581 247 249 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
* Pins of element D2580 are shorted:
* D2580 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -778 -1605.499 -774)CMOSN2580 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2579 are shorted:
* D2579 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -762 -1605.499 -758)CMOSN2579 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2578 are shorted:
* D2578 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -746 -1605.499 -742)CMOSN2578 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2577 are shorted:
* D2577 8 8 D_lateral AREA=8.625f    ; (-1668.5 -730 -1605.499 -718)CMOSN2577 8 8 D_lateral AREA=8.625f    
* Pins of element D2576 are shorted:
* D2576 8 8 D_lateral AREA=4.375E-016    ; (-1673.501 -726 -1673.5 -719)CMOSN2576 8 8 D_lateral AREA=4.375E-016    
* Pins of element D2575 are shorted:
* D2575 8 8 D_lateral AREA=4.1250625f    ; (-1673.501 -706 -1615.5 -697.999)CMOSN2575 8 8 D_lateral AREA=4.1250625f    
M2574 248 247 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M2573 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2572 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2571 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2570 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2569 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2568 248 247 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M2567 247 249 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M2566 247 249 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D2565 are shorted:
* D2565 12 12 D_lateral AREA=2.4374375f    ; (-1730.5 -706 -1697.5 -700)CMOSN2565 12 12 D_lateral AREA=2.4374375f    
* Pins of element D2564 are shorted:
* D2564 12 12 D_lateral AREA=2.687375f    ; (-1732.5 -722 -1697.5 -718)CMOSN2564 12 12 D_lateral AREA=2.687375f    
* Pins of element D2563 are shorted:
* D2563 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -778 -1733.499 -774)CMOSN2563 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2562 are shorted:
* D2562 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -762 -1733.499 -758)CMOSN2562 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2561 are shorted:
* D2561 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -746 -1733.499 -742)CMOSN2561 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2560 are shorted:
* D2560 12 12 D_lateral AREA=2.3749375f    ; (-1733.5 -730 -1699.5 -726)CMOSN2560 12 12 D_lateral AREA=2.3749375f    
C2557 249 12  184.041f    ; (-2185.5 -787 -1899.5 -501)CMOSN.041f    
M2556 8 389 404 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2555 256 250 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2554 389 390 256 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2553 255 399 390 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2552 8 401 255 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2550 8 262 254 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2549 254 260 250 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2547 389 250 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2546 12 390 389 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2545 12 262 250 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2544 250 260 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2542 12 251 267 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2541 12 264 252 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2540 252 253 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2538 8 285 399 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2537 8 285 257 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2536 257 402 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2535 8 402 401 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2534 257 401 403 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2533 257 399 403 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2532 8 267 260 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2531 8 267 259 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2530 259 268 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2529 8 268 262 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2528 259 262 402 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2527 259 260 402 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2526 12 267 260 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2525 258 267 402 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2524 258 268 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2523 12 268 262 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2522 258 262 402 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2521 12 260 258 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2520 12 172 253 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2519 261 172 265 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2518 261 263 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2517 12 263 264 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2516 261 264 265 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2515 12 253 261 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2514 8 269 268 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2511 8 73 165 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2510 165 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2509 408 410 271 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2507 12 269 268 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2505 270 248 165 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2504 12 73 270 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2503 12 410 408 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
* Pins of element D2501 are shorted:
* D2501 12 12 D_lateral AREA=3.125E-016    ; (696.5 -823 701.5 -822.999)CMOSN2501 12 12 D_lateral AREA=3.125E-016    
M2500 8 408 425 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2499 8 273 271 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=562.5f PS=2.25u    
M2498 277 419 410 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2497 8 422 277 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2496 419 310 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2495 8 310 278 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2494 8 282 276 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2493 276 289 273 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2492 289 288 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2491 8 288 280 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2490 12 273 408 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=968.75f PS=3u    
M2489 12 282 273 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2488 273 289 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2487 289 288 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2486 12 289 279 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2485 12 272 288 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2484 12 284 274 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2483 274 275 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2482 275 188 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2481 12 275 281 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2480 8 429 292 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2479 278 423 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2478 8 423 422 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2477 278 422 420 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2476 278 419 420 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2475 280 292 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2474 8 292 282 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2473 280 282 423 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2472 280 289 423 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2471 12 429 292 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2469 279 292 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2468 12 292 282 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2467 279 282 423 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2466 279 288 423 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2465 287 248 290 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2464 12 83 287 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2463 281 283 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2462 12 283 284 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2461 281 284 285 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2460 281 188 285 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D2459 are shorted:
* D2459 12 12 D_lateral AREA=3.125E-016    ; (412 -823 417 -822.999)CMOSN2459 12 12 D_lateral AREA=3.125E-016    
M2456 8 83 290 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2455 290 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2454 8 430 445 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2453 293 296 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2452 430 434 293 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2451 430 296 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2450 12 434 430 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2449 12 291 295 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2448 300 432 434 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2447 8 440 300 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2446 432 329 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2445 8 329 301 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2444 301 432 427 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2443 8 306 299 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2442 299 294 296 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2441 294 295 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2440 8 295 303 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2439 303 294 441 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2438 12 306 296 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2437 296 294 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2436 294 295 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2435 302 295 441 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2434 12 294 302 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2433 12 309 297 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2432 297 298 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2431 298 192 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2430 304 192 310 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2429 12 298 304 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2428 8 439 305 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2427 301 441 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2426 8 441 440 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2425 301 440 427 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2424 303 305 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2423 8 305 306 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2422 303 306 441 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2421 12 439 305 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2419 302 305 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2418 12 305 306 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2417 302 306 441 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2416 312 248 307 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2415 12 18 312 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2414 304 308 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2413 12 308 309 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2412 304 309 310 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
* Pins of element D2411 are shorted:
* D2411 12 12 D_lateral AREA=3.125E-016    ; (128 -823 133 -822.999)CMOSN2411 12 12 D_lateral AREA=3.125E-016    
M2408 8 18 307 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2407 307 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2406 8 452 457 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2405 314 321 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2404 452 459 314 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2403 452 321 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2402 12 459 452 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2401 12 313 320 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2400 326 455 459 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2399 8 466 326 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2398 455 354 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2397 8 354 315 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2396 315 466 467 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2394 315 455 467 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2393 8 327 325 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2392 325 316 321 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2391 316 320 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2390 8 320 318 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2389 318 327 469 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2387 318 316 469 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2386 12 327 321 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2385 321 316 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2384 316 320 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2383 317 320 469 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2382 317 327 469 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2380 12 316 317 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2379 12 332 322 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2378 322 324 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2377 324 220 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2376 319 220 329 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2375 319 332 329 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2373 12 324 319 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2372 8 468 328 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2371 8 469 315 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2370 8 469 466 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2369 8 328 318 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2368 8 328 327 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2367 12 468 328 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2365 12 328 317 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2364 12 328 327 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2363 333 248 330 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2362 12 334 333 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2361 12 331 319 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M2360 12 331 332 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D2359 are shorted:
* D2359 12 12 D_lateral AREA=3.125E-016    ; (-156.5 -823 -151.5 -822.999)CMOSN2359 12 12 D_lateral AREA=3.125E-016    
M2356 8 334 330 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2355 330 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2354 8 473 481 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2353 338 345 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2352 473 483 338 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2350 8 487 337 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2349 8 349 336 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2347 473 345 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2346 12 483 473 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2345 12 349 345 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2344 12 335 344 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2343 12 350 346 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2342 483 479 337 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2341 479 373 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2340 8 373 339 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2339 339 487 490 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2338 339 489 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2337 8 489 487 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2336 339 479 490 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2335 345 340 336 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2334 340 344 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2333 8 344 342 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2332 342 349 489 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2331 342 351 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2330 8 351 349 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2329 342 340 489 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2328 345 340 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2327 340 344 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2326 341 344 489 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2325 341 349 489 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2324 341 351 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2323 12 351 349 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2322 12 340 341 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2321 346 348 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2320 348 228 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2319 343 228 354 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2318 343 350 354 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2317 343 353 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2316 12 353 350 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2315 12 348 343 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2314 8 488 351 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2312 8 37 352 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2311 12 488 351 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2309 355 248 352 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2308 12 37 355 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2307 are shorted:
* D2307 12 12 D_lateral AREA=3.125E-016    ; (-441 -823 -436 -822.999)CMOSN2307 12 12 D_lateral AREA=3.125E-016    
M2305 352 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2304 8 494 507 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2303 361 356 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2302 494 495 361 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2301 360 505 495 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2300 8 509 360 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2299 8 368 359 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2298 359 363 356 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2297 494 356 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2296 12 495 494 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2295 12 368 356 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2294 356 363 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2293 12 357 367 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2292 12 369 358 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2291 358 371 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2290 505 381 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2289 8 381 362 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2288 362 374 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2287 8 374 509 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2286 362 509 511 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2285 362 505 511 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2284 363 367 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2283 8 367 365 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2282 365 372 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2281 8 372 368 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2280 365 368 374 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2279 365 363 374 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2278 363 367 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2277 364 367 374 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2276 364 372 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2275 12 372 368 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2274 364 368 374 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2273 12 363 364 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2272 371 238 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2271 366 238 373 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2270 366 236 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2269 12 236 369 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2268 366 369 373 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2267 12 371 366 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2266 8 512 372 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2263 8 40 375 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2262 375 248 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2261 12 512 372 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2259 376 248 375 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2258 12 40 376 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2257 are shorted:
* D2257 12 12 D_lateral AREA=3.125E-016    ; (-725.5 -823 -720.5 -822.999)CMOSN2257 12 12 D_lateral AREA=3.125E-016    
M2256 8 382 377 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2255 377 380 516 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2254 12 382 516 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2253 516 380 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2252 380 383 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2251 8 383 379 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2250 379 384 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2249 8 384 382 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2248 379 382 522 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2247 379 380 522 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2246 380 383 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2245 378 383 522 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2244 378 384 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2243 12 384 382 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2242 378 382 522 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2241 12 380 378 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2240 8 41 384 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2239 384 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2238 385 442 384 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2237 12 41 385 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2236 are shorted:
* D2236 12 12 D_lateral AREA=3.125E-016    ; (-1002.5 -894 -997.5 -893.999)CMOSN2236 12 12 D_lateral AREA=3.125E-016    
M2224 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2223 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2222 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2221 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2220 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2219 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M2218 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D2217 are shorted:
* D2217 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1000 1697.5 -996)CMOSN2217 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2216 are shorted:
* D2216 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -984 1697.5 -980)CMOSN2216 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2215 are shorted:
* D2215 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -968 1697.5 -964)CMOSN2215 12 12 D_lateral AREA=2.5E-016    
* Pins of element D2214 are shorted:
* D2214 12 12 D_lateral AREA=3.249875f    ; (1661.5 -952 1697.5 -944)CMOSN2214 12 12 D_lateral AREA=3.249875f    
* Pins of element D2213 are shorted:
* D2213 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -997 1637.501 -993)CMOSN2213 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2212 are shorted:
* D2212 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -981 1637.501 -977)CMOSN2212 8 8 D_lateral AREA=2.5E-016    
* Pins of element D2211 are shorted:
* D2211 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -965 1637.501 -961)CMOSN2211 8 8 D_lateral AREA=2.5E-016    
M2209 386 387 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M2207 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2205 386 387 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M2203 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2201 386 387 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M2199 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2197 386 387 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M2194 386 387 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M2193 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2192 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2191 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2190 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2189 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M2188 8 387 386 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D2187 are shorted:
* D2187 8 8 D_lateral AREA=8.875125f    ; (1502.499 -949 1637.501 -944.999)CMOSN2187 8 8 D_lateral AREA=8.875125f    
M2186 8 530 541 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2185 393 388 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2184 530 528 393 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2183 392 529 528 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2182 8 540 392 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2181 8 400 391 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2180 391 397 388 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2179 530 388 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2178 12 528 530 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2177 12 400 388 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2176 388 397 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2175 12 389 404 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2174 12 401 390 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2173 390 399 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2171 529 420 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2170 8 420 394 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2169 394 539 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2168 8 539 540 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2167 394 540 537 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2166 394 529 537 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2165 397 404 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2164 8 404 396 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2163 396 405 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2162 8 405 400 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2161 396 400 539 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2160 396 397 539 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2159 397 404 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2158 395 404 539 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2157 395 405 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2156 12 405 400 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2155 395 400 539 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2154 12 397 395 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2153 12 285 399 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2152 398 285 403 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2151 398 402 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2150 12 402 401 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2149 398 401 403 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2148 12 399 398 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2147 8 73 405 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2146 405 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2145 8 73 269 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2144 269 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2143 407 696 405 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2142 12 73 407 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2140 406 442 269 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2139 12 73 406 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D2138 are shorted:
* D2138 12 12 D_lateral AREA=3.125E-016    ; (696.5 -964 701.5 -963.999)CMOSN2138 12 12 D_lateral AREA=3.125E-016    
* Pins of element D2137 are shorted:
* D2137 12 12 D_lateral AREA=3.125E-016    ; (696.5 -919 701.5 -918.999)CMOSN2137 12 12 D_lateral AREA=3.125E-016    
M2136 8 545 558 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2135 413 409 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2134 545 543 413 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2133 412 544 543 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2132 8 557 412 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2131 8 427 544 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2130 8 421 411 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2129 411 417 409 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2128 8 425 417 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M2127 545 409 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2126 545 543 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.9375p PS=6u    
M2125 12 421 409 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2124 409 417 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2123 12 425 417 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M2122 12 408 425 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2121 12 422 410 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2120 410 419 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2119 419 310 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2118 12 419 418 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2117 414 556 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2116 8 556 557 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2115 414 557 554 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2114 414 544 554 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2113 8 427 414 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2112 416 428 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2111 8 428 421 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2110 416 421 556 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2109 416 417 556 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2108 8 425 416 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2107 426 696 428 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2106 12 83 426 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2105 415 428 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2104 12 428 421 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2103 415 421 556 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2102 12 417 415 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2101 415 425 556 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2100 424 442 429 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2099 12 83 424 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2098 418 423 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2097 12 423 422 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2096 418 422 420 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2095 418 310 420 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
* Pins of element D2094 are shorted:
* D2094 12 12 D_lateral AREA=3.125E-016    ; (412 -964 417 -963.999)CMOSN2094 12 12 D_lateral AREA=3.125E-016    
* Pins of element D2093 are shorted:
* D2093 12 12 D_lateral AREA=3.125E-016    ; (412 -919 417 -918.999)CMOSN2093 12 12 D_lateral AREA=3.125E-016    
M2092 8 560 573 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2091 431 433 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2090 560 563 431 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2089 8 83 428 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2088 428 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2087 8 83 429 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2086 429 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2085 560 433 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2084 12 563 560 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2083 12 430 445 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2082 436 450 563 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2081 8 571 436 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2080 450 467 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2079 8 467 449 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2078 8 438 435 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2077 435 448 433 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2076 448 445 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2075 8 445 447 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2074 12 438 433 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2073 433 448 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2072 448 445 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2071 12 448 444 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2070 12 440 434 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2069 434 432 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2068 432 329 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2067 437 329 427 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2066 12 432 437 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2065 449 569 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2064 8 569 571 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2063 449 571 566 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2062 449 450 566 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2061 447 451 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2060 8 451 438 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2059 447 438 569 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2058 447 448 569 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2057 446 696 451 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2056 12 18 446 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2055 444 451 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2054 12 451 438 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2053 444 438 569 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2052 444 445 569 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2051 443 442 439 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2050 12 18 443 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2049 437 441 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2048 12 441 440 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2047 437 440 427 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
* Pins of element D2046 are shorted:
* D2046 12 12 D_lateral AREA=3.125E-016    ; (128 -964 133 -963.999)CMOSN2046 12 12 D_lateral AREA=3.125E-016    
* Pins of element D2045 are shorted:
* D2045 12 12 D_lateral AREA=3.125E-016    ; (128 -919 133 -918.999)CMOSN2045 12 12 D_lateral AREA=3.125E-016    
M2044 8 577 580 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M2043 453 458 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M2042 577 581 453 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M2041 8 18 451 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2040 451 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2039 8 18 439 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M2038 439 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M2037 577 458 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M2036 12 581 577 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M2035 12 452 457 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M2034 461 584 581 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2033 8 582 461 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2032 584 490 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2031 8 490 462 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2029 462 584 592 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2028 8 463 460 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M2027 460 454 458 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M2026 454 457 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M2025 8 457 465 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M2023 465 454 594 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M2022 12 463 458 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2021 458 454 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2020 454 457 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2019 464 457 594 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2017 12 454 464 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2016 12 466 459 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M2015 459 455 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M2014 455 354 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M2013 456 354 467 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M2012 456 466 467 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M2010 12 455 456 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M2009 462 594 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2008 8 594 582 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2007 462 582 592 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2006 465 472 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2005 8 472 463 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M2004 465 463 594 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M2003 471 696 472 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M2002 12 334 471 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M2001 464 472 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M2000 12 472 463 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1999 464 463 594 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1998 470 442 468 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1997 12 334 470 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1996 12 469 456 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=968.75f PS=3u    
M1995 12 469 466 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
* Pins of element D1994 are shorted:
* D1994 12 12 D_lateral AREA=3.125E-016    ; (-156.5 -964 -151.5 -963.999)CMOSN1994 12 12 D_lateral AREA=3.125E-016    
* Pins of element D1993 are shorted:
* D1993 12 12 D_lateral AREA=3.125E-016    ; (-156.5 -919 -151.5 -918.999)CMOSN1993 12 12 D_lateral AREA=3.125E-016    
M1992 8 595 602 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1991 474 482 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1990 595 603 474 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1989 8 334 472 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1988 472 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1987 8 334 468 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1986 468 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1985 595 482 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1984 12 603 595 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1983 12 473 481 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1982 12 487 483 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1981 485 606 603 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1980 8 605 485 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1979 606 511 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1978 8 511 475 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1977 475 605 610 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1976 475 612 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1975 475 606 610 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1974 8 486 484 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1973 484 476 482 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1972 476 481 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1971 8 481 478 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1970 478 486 612 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1969 478 493 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1968 478 476 612 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1967 12 486 482 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1966 482 476 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1965 476 481 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1964 477 481 612 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1963 477 486 612 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1962 477 493 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1961 12 476 477 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1960 483 479 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1959 479 373 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1958 480 373 490 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1957 480 487 490 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1956 480 489 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1955 12 489 487 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1954 12 479 480 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1953 8 37 493 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1952 8 612 605 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1951 8 493 486 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1950 8 37 488 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1949 492 696 493 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1948 12 37 492 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1947 12 493 486 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1946 491 442 488 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1945 12 37 491 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1944 are shorted:
* D1944 12 12 D_lateral AREA=3.125E-016    ; (-441 -964 -436 -963.999)CMOSN1944 12 12 D_lateral AREA=3.125E-016    
* Pins of element D1943 are shorted:
* D1943 12 12 D_lateral AREA=3.125E-016    ; (-441 -919 -436 -918.999)CMOSN1943 12 12 D_lateral AREA=3.125E-016    
M1942 8 613 624 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1941 498 502 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1940 613 499 498 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1939 497 626 499 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1938 8 627 497 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1937 8 508 496 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1936 496 501 502 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1935 493 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1934 488 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1933 613 502 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1932 12 499 613 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1931 12 508 502 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1929 12 494 507 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1928 12 509 495 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1927 495 505 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1926 626 522 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1925 8 522 500 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1924 500 627 628 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1923 500 629 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1922 8 629 627 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1921 500 626 628 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1920 501 507 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1919 8 507 504 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1918 504 508 629 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1917 504 510 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1916 8 510 508 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1915 504 501 629 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1914 12 501 502 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1913 501 507 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1912 503 507 629 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1911 503 508 629 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1910 503 510 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1909 12 510 508 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1908 12 501 503 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1907 505 381 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1906 506 381 511 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1905 506 374 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1904 12 374 509 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1903 506 509 511 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1902 12 505 506 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1901 8 40 510 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1900 510 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1899 8 40 512 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1898 512 442 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1897 514 696 510 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1896 12 40 514 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
M1895 513 442 512 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1894 12 40 513 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1893 are shorted:
* D1893 12 12 D_lateral AREA=3.125E-016    ; (-725.5 -964 -720.5 -963.999)CMOSN1893 12 12 D_lateral AREA=3.125E-016    
* Pins of element D1892 are shorted:
* D1892 12 12 D_lateral AREA=3.125E-016    ; (-725.5 -919 -720.5 -918.999)CMOSN1892 12 12 D_lateral AREA=3.125E-016    
M1891 8 523 517 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1890 517 515 682 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1889 515 516 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1888 8 516 519 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1887 519 515 521 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1886 12 523 682 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1885 682 515 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1884 515 516 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1883 518 516 521 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1882 12 515 518 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1881 519 520 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1880 8 520 523 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1879 519 523 521 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1878 520 524 8 8 CMOSP L=750n W=2.25u AD=2.46875p PD=7.25u AS=2.46875p PS=7.25u    
M1877 518 520 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1876 12 520 523 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1875 518 523 521 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1874 520 524 12 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=1.75p PS=5.5u    
M1873 8 41 524 8 CMOSP L=1.25u W=5u AD=7.5p PD=13u AS=5.625p PS=7.25u    
M1872 524 696 8 8 CMOSP L=1.25u W=5u AD=5.625p PD=7.25u AS=7.5p PS=13u    
M1871 525 696 524 12 CMOSN L=1.25u W=1.25u AD=468.75f PD=2u AS=2.65625p PS=6.75u    
M1870 12 41 525 12 CMOSN L=1.25u W=1.25u AD=1.5625p PD=5u AS=468.75f PS=2u    
* Pins of element D1869 are shorted:
* D1869 12 12 D_lateral AREA=3.125E-016    ; (-1002.5 -989 -997.5 -988.999)CMOSN1869 12 12 D_lateral AREA=3.125E-016    
M1859 8 526 684 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1857 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1855 8 526 684 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1853 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1851 8 526 684 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1849 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1847 8 526 684 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1845 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1842 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M1841 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1840 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1839 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1838 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1837 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1836 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1835 684 526 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1833 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1832 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1831 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1830 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1829 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1828 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1827 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D1826 are shorted:
* D1826 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -996 -1760.499 -992)CMOSN1826 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1825 are shorted:
* D1825 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -980 -1760.499 -976)CMOSN1825 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1824 are shorted:
* D1824 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -964 -1760.499 -960)CMOSN1824 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1823 are shorted:
* D1823 12 12 D_lateral AREA=3.249875f    ; (-1760.5 -948 -1724.5 -940)CMOSN1823 12 12 D_lateral AREA=3.249875f    
* Pins of element D1821 are shorted:
* D1821 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -993 -1700.5 -989)CMOSN1821 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1820 are shorted:
* D1820 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -977 -1700.5 -973)CMOSN1820 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1819 are shorted:
* D1819 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -961 -1700.5 -957)CMOSN1819 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1818 are shorted:
* D1818 8 8 D_lateral AREA=8.875125f    ; (-1700.501 -945 -1565.499 -940.999)CMOSN1818 8 8 D_lateral AREA=8.875125f    
M1809 387 8 643 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M1808 643 8 387 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M1807 387 8 643 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M1806 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1805 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1804 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1803 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1802 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1801 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1800 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1799 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1798 386 643 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1797 643 265 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1796 12 265 643 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1795 643 265 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M1794 12 527 643 12 CMOSN L=500n W=3u AD=6.0625p PD=10.75u AS=2.25p PS=4.5u    
* Pins of element D1792 are shorted:
* D1792 12 12 D_lateral AREA=2.3749375f    ; (1663.5 -1080 1697.5 -1076)CMOSN1792 12 12 D_lateral AREA=2.3749375f    
* Pins of element D1791 are shorted:
* D1791 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1064 1697.5 -1060)CMOSN1791 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1790 are shorted:
* D1790 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1048 1697.5 -1044)CMOSN1790 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1789 are shorted:
* D1789 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1032 1697.5 -1028)CMOSN1789 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1788 are shorted:
* D1788 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1016 1697.5 -1012)CMOSN1788 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1787 are shorted:
* D1787 8 8 D_lateral AREA=1.8125625f    ; (1614.5 -1015.001 1637.501 -1009)CMOSN1787 8 8 D_lateral AREA=1.8125625f    
* Pins of element D1786 are shorted:
* D1786 8 8 D_lateral AREA=3.125E-016    ; (1611.5 -1073 1611.501 -1068)CMOSN1786 8 8 D_lateral AREA=3.125E-016    
M1785 387 265 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M1784 387 265 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M1783 387 265 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M1782 643 527 387 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M1781 387 527 643 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M1780 643 527 387 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M1779 387 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M1778 8 387 386 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
* Pins of element D1776 are shorted:
* D1776 8 8 D_lateral AREA=3.125E-016    ; (1558.499 -1073 1558.5 -1068)CMOSN1776 8 8 D_lateral AREA=3.125E-016    
* Pins of element D1775 are shorted:
* D1775 8 8 D_lateral AREA=2.5E-016    ; (1558.499 -1056 1558.5 -1052)CMOSN1775 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1774 are shorted:
* D1774 8 8 D_lateral AREA=3.5625625f    ; (1558.499 -1040 1605.5 -1029.999)CMOSN1774 8 8 D_lateral AREA=3.5625625f    
M1773 8 387 386 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1772 8 538 531 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1771 531 535 559 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1770 12 530 541 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1769 12 540 528 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1768 528 529 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1767 12 538 559 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1766 559 535 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1765 535 541 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1764 8 541 534 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1763 534 554 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1762 8 554 538 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1761 534 538 536 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1760 534 535 536 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1759 532 540 537 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1758 12 539 540 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1757 529 420 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1756 532 420 537 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1755 12 529 532 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1754 532 539 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1753 535 541 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1752 533 541 536 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1751 533 554 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1750 12 554 538 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1749 533 538 536 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1748 12 535 533 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1746 8 645 568 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1745 548 542 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1744 645 646 548 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1743 547 648 646 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1742 8 649 547 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1741 8 559 648 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M1740 8 555 546 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1739 546 552 542 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1738 8 558 552 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=2.21875p PS=6.75u    
M1737 645 542 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1736 645 646 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.9375p PS=6u    
M1735 12 555 542 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1734 542 552 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1733 12 558 552 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=2.21875p PS=6.75u    
M1732 12 545 558 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1731 12 557 543 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1730 543 544 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1729 544 427 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1728 549 650 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1727 8 650 649 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1726 549 649 698 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1725 549 648 698 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1724 8 559 549 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1723 551 566 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1722 8 566 555 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1721 551 555 650 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1720 551 552 650 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1719 8 558 551 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1718 550 566 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1717 12 566 555 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1716 550 555 650 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1715 12 552 550 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1714 550 558 650 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1713 553 557 554 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1712 12 556 557 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1711 553 427 554 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1710 12 544 553 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1709 553 556 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1708 8 651 593 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1707 561 562 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1706 651 652 561 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1705 651 562 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1704 12 652 651 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1703 12 560 573 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1702 565 653 652 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1701 8 654 565 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1700 653 568 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1699 8 568 576 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1698 8 567 564 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1697 564 575 562 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1696 575 573 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1695 8 573 574 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1694 12 567 562 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1693 562 575 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1692 575 573 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1691 12 575 572 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1690 12 571 563 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1689 563 450 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1688 450 467 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1687 12 450 570 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1686 576 655 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1685 8 655 654 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1684 576 654 699 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1683 576 653 699 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1682 574 592 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1681 8 592 567 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1680 574 567 655 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1679 574 575 655 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1678 572 592 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1677 12 592 567 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1676 572 567 655 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1675 572 573 655 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1674 570 571 566 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1673 12 569 571 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1672 570 467 566 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1671 570 569 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1670 8 657 611 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1669 578 583 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1668 657 659 578 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1667 12 577 580 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1666 657 583 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1665 12 659 657 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1664 586 658 659 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1663 8 660 586 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1662 658 593 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1661 8 593 588 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1659 588 658 687 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1658 8 589 585 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1657 585 579 583 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1656 579 580 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1655 8 580 591 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1653 591 579 662 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1652 12 582 581 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1651 581 584 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1649 584 490 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1648 587 490 592 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1647 12 584 587 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1646 12 589 583 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1645 583 579 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1644 579 580 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1643 590 580 662 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1641 12 579 590 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1640 588 662 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1639 8 662 660 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1638 588 660 687 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1637 591 610 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1636 8 610 589 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1635 591 589 662 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1634 587 582 592 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1633 12 594 582 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1632 587 594 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1631 590 610 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1630 12 610 589 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1629 590 589 662 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1628 8 663 673 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1627 596 604 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1626 663 666 596 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1625 12 595 602 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1624 663 604 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1623 12 666 663 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1622 608 664 666 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1621 8 667 608 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1620 664 611 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1619 8 611 598 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1618 598 667 734 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1617 598 668 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1616 598 664 734 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1615 8 609 607 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1614 607 599 604 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1613 599 602 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1612 8 602 601 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1611 601 609 668 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1610 601 628 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1609 601 599 668 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1608 12 605 603 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1607 603 606 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1606 597 605 610 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1605 606 511 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1604 597 511 610 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1603 12 606 597 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1602 597 612 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1601 12 609 604 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1600 604 599 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1599 599 602 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1598 600 602 668 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1597 600 609 668 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1596 600 628 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1595 12 599 600 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1594 8 668 667 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1593 8 628 609 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1592 12 612 605 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1591 12 628 609 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1590 8 669 639 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1589 616 621 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1588 669 618 616 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1587 615 670 618 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1586 8 672 615 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1585 8 625 614 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1584 614 620 621 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1583 12 613 624 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1582 12 627 499 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1580 669 621 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1579 12 618 669 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1578 12 625 621 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1576 670 673 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1575 8 673 619 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1574 619 672 741 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1573 619 674 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1572 8 674 672 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1571 619 670 741 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1570 620 624 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1569 8 624 623 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1568 623 625 674 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1567 623 521 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1566 8 521 625 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1565 623 620 674 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1564 12 626 499 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1563 617 627 628 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1562 12 629 627 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1561 626 522 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1560 617 522 628 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1559 12 626 617 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1558 617 629 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1557 12 620 621 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1556 620 624 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1555 622 624 674 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1554 622 625 674 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1553 622 521 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1552 12 521 625 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1551 12 620 622 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1550 8 675 676 8 CMOSP L=750n W=1.5u AD=2.25p PD=6u AS=2.25p PS=6u    
M1549 633 630 8 8 CMOSP L=750n W=750n AD=562.5f PD=2.25u AS=1.75p PS=5.5u    
M1548 675 677 633 8 CMOSP L=750n W=750n AD=2.3125p PD=7u AS=562.5f PS=2.25u    
M1547 632 679 677 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1546 8 680 632 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1545 8 638 631 8 CMOSP L=750n W=750n AD=1.75p PD=5.5u AS=187.5f PS=1.25u    
M1544 631 637 630 8 CMOSP L=750n W=750n AD=187.5f PD=1.25u AS=1.75p PS=5.5u    
M1543 675 630 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.90625p PS=5.75u    
M1542 12 677 675 12 CMOSN L=750n W=750n AD=1.9375p PD=6u AS=968.75f PS=3u    
M1541 12 638 630 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1540 630 637 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1539 679 682 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1538 8 682 634 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1537 634 681 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1536 8 681 680 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1535 634 680 747 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1534 634 679 747 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1533 637 639 8 8 CMOSP L=750n W=750n AD=2.21875p PD=6.75u AS=1.15625p PS=3.5u    
M1532 8 639 636 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.109375p PS=3.375u    
M1531 636 8 8 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1530 8 8 638 8 CMOSP L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1529 636 638 681 8 CMOSP L=750n W=750n AD=968.75f PD=3u AS=7.4375p PS=19.125u    
M1528 636 637 681 8 CMOSP L=750n W=750n AD=1.109375p PD=3.375u AS=7.4375p PS=19.125u    
M1527 637 639 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1526 635 639 681 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1525 635 8 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1524 12 8 638 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1523 635 638 681 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1522 12 637 635 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1521 8 12 526 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M1520 526 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M1519 526 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M1518 640 641 526 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M1517 526 641 640 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M1516 640 641 526 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M1515 526 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
* Pins of element D1513 are shorted:
* D1513 8 8 D_lateral AREA=2.5E-016    ; (-1621.5 -1052 -1621.499 -1048)CMOSN1513 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1512 are shorted:
* D1512 8 8 D_lateral AREA=3.5625625f    ; (-1668.5 -1036 -1621.499 -1025.999)CMOSN1512 8 8 D_lateral AREA=3.5625625f    
* Pins of element D1511 are shorted:
* D1511 8 8 D_lateral AREA=3.125E-016    ; (-1621.5 -1069 -1621.499 -1064)CMOSN1511 8 8 D_lateral AREA=3.125E-016    
* Pins of element D1510 are shorted:
* D1510 8 8 D_lateral AREA=3.125E-016    ; (-1674.501 -1069 -1674.5 -1064)CMOSN1510 8 8 D_lateral AREA=3.125E-016    
M1509 640 12 526 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M1508 526 12 640 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M1507 640 12 526 12 CMOSN L=500n W=3.25u AD=2.53125p PD=5u AS=4.875p PS=9.5u    
M1506 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1505 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1504 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1503 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1502 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1501 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1500 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1499 684 640 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1498 12 640 684 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1497 640 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1496 12 12 640 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1495 640 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M1494 640 641 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D1491 are shorted:
* D1491 12 12 D_lateral AREA=2.3749375f    ; (-1760.5 -1076 -1726.5 -1072)CMOSN1491 12 12 D_lateral AREA=2.3749375f    
* Pins of element D1490 are shorted:
* D1490 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1060 -1760.499 -1056)CMOSN1490 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1489 are shorted:
* D1489 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1044 -1760.499 -1040)CMOSN1489 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1488 are shorted:
* D1488 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1028 -1760.499 -1024)CMOSN1488 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1487 are shorted:
* D1487 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1012 -1760.499 -1008)CMOSN1487 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1486 are shorted:
* D1486 8 8 D_lateral AREA=1.8125625f    ; (-1700.501 -1011.001 -1677.5 -1005)CMOSN1486 8 8 D_lateral AREA=1.8125625f    
M1478 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1477 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1476 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1475 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1474 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1473 527 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M1472 642 386 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M1471 642 386 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D1470 are shorted:
* D1470 12 12 D_lateral AREA=3.75E-016    ; (1632.5 -1112 1632.501 -1106)CMOSN1470 12 12 D_lateral AREA=3.75E-016    
* Pins of element D1469 are shorted:
* D1469 12 12 D_lateral AREA=2f    ; (1641.499 -1115 1651.5 -1103)CMOSN1469 12 12 D_lateral AREA=2f    
* Pins of element D1468 are shorted:
* D1468 12 12 D_lateral AREA=2.687375f    ; (1634.5 -1162 1669.5 -1158)CMOSN1468 12 12 D_lateral AREA=2.687375f    
* Pins of element D1467 are shorted:
* D1467 12 12 D_lateral AREA=2.4374375f    ; (1634.5 -1146 1667.5 -1140)CMOSN1467 12 12 D_lateral AREA=2.4374375f    
* Pins of element D1466 are shorted:
* D1466 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1202 1670.5 -1198)CMOSN1466 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1465 are shorted:
* D1465 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1186 1670.5 -1182)CMOSN1465 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1464 are shorted:
* D1464 12 12 D_lateral AREA=2.3749375f    ; (1636.5 -1170 1670.5 -1166)CMOSN1464 12 12 D_lateral AREA=2.3749375f    
M1462 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1461 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1460 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1459 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1458 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1457 642 386 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1456 642 386 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M1455 527 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D1454 are shorted:
* D1454 8 8 D_lateral AREA=4.1250625f    ; (1552.5 -1146 1610.501 -1137.999)CMOSN1454 8 8 D_lateral AREA=4.1250625f    
* Pins of element D1453 are shorted:
* D1453 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1202 1542.5 -1198)CMOSN1453 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1452 are shorted:
* D1452 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1186 1542.5 -1182)CMOSN1452 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1451 are shorted:
* D1451 8 8 D_lateral AREA=4.375E-016    ; (1610.5 -1166 1610.501 -1159)CMOSN1451 8 8 D_lateral AREA=4.375E-016    
* Pins of element D1450 are shorted:
* D1450 8 8 D_lateral AREA=8.625f    ; (1542.499 -1170 1605.5 -1158)CMOSN1450 8 8 D_lateral AREA=8.625f    
* Pins of element D1449 are shorted:
* D1449 8 8 D_lateral AREA=4.062625f    ; (1558.499 -1128.001 1611.501 -1122)CMOSN1449 8 8 D_lateral AREA=4.062625f    
M1448 12 645 568 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1447 12 649 646 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1446 646 648 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1445 648 559 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1444 647 649 698 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1443 12 650 649 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1442 12 648 647 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1441 647 559 698 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1440 647 650 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1439 12 651 593 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1438 12 654 652 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1437 652 653 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1436 12 653 656 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1435 653 568 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1434 656 654 699 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1433 12 655 654 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1432 656 568 699 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1431 656 655 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1430 12 657 611 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1429 12 660 659 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1428 659 658 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1426 12 658 661 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1425 658 593 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1424 661 593 687 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1423 661 660 687 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1422 12 662 660 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1421 661 662 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1420 12 663 673 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1419 12 667 666 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1418 666 664 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1417 665 667 734 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1416 12 664 665 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1415 664 611 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1414 665 611 734 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1413 665 668 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1412 12 668 667 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1411 12 669 639 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1410 12 672 618 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1408 12 670 618 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1407 671 672 741 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1406 12 674 672 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1405 12 670 671 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1404 670 673 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1403 671 673 741 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1402 671 674 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1401 12 675 676 12 CMOSN L=750n W=750n AD=1.90625p PD=5.75u AS=1.75p PS=5.5u    
M1400 12 680 677 12 CMOSN L=750n W=750n AD=1.75p PD=5.5u AS=968.75f PS=3u    
M1399 677 679 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.75p PS=5.5u    
M1398 678 680 747 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=7.375p PS=19u    
M1397 12 681 680 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=1.75p PS=5.5u    
M1396 12 679 678 12 CMOSN L=750n W=750n AD=1.109375p PD=3.375u AS=1.15625p PS=3.5u    
M1395 679 682 12 12 CMOSN L=750n W=750n AD=2.21875p PD=6.75u AS=1.109375p PS=3.375u    
M1394 678 682 747 12 CMOSN L=750n W=750n AD=1.15625p PD=3.5u AS=7.375p PS=19u    
M1393 678 681 12 12 CMOSN L=750n W=750n AD=968.75f PD=3u AS=1.15625p PS=3.5u    
M1392 442 683 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1391 8 683 442 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M1390 442 683 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1389 8 683 442 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M1388 442 683 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1387 683 684 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1386 683 684 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M1385 641 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D1384 are shorted:
* D1384 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1198 -1605.499 -1194)CMOSN1384 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1383 are shorted:
* D1383 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1182 -1605.499 -1178)CMOSN1383 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1382 are shorted:
* D1382 8 8 D_lateral AREA=8.625f    ; (-1668.5 -1166 -1605.499 -1154)CMOSN1382 8 8 D_lateral AREA=8.625f    
* Pins of element D1381 are shorted:
* D1381 8 8 D_lateral AREA=4.375E-016    ; (-1673.501 -1162 -1673.5 -1155)CMOSN1381 8 8 D_lateral AREA=4.375E-016    
* Pins of element D1380 are shorted:
* D1380 8 8 D_lateral AREA=4.1250625f    ; (-1673.501 -1142 -1615.5 -1133.999)CMOSN1380 8 8 D_lateral AREA=4.1250625f    
* Pins of element D1379 are shorted:
* D1379 8 8 D_lateral AREA=4.062625f    ; (-1674.501 -1124.001 -1621.499 -1118)CMOSN1379 8 8 D_lateral AREA=4.062625f    
M1378 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1377 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1376 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1375 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1374 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1373 641 12 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M1372 683 684 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M1371 683 684 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D1370 are shorted:
* D1370 12 12 D_lateral AREA=3.75E-016    ; (-1695.501 -1108 -1695.5 -1102)CMOSN1370 12 12 D_lateral AREA=3.75E-016    
* Pins of element D1369 are shorted:
* D1369 12 12 D_lateral AREA=2f    ; (-1714.5 -1111 -1704.499 -1099)CMOSN1369 12 12 D_lateral AREA=2f    
* Pins of element D1368 are shorted:
* D1368 12 12 D_lateral AREA=2.4374375f    ; (-1730.5 -1142 -1697.5 -1136)CMOSN1368 12 12 D_lateral AREA=2.4374375f    
* Pins of element D1367 are shorted:
* D1367 12 12 D_lateral AREA=2.687375f    ; (-1732.5 -1158 -1697.5 -1154)CMOSN1367 12 12 D_lateral AREA=2.687375f    
* Pins of element D1366 are shorted:
* D1366 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1198 -1733.499 -1194)CMOSN1366 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1365 are shorted:
* D1365 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1182 -1733.499 -1178)CMOSN1365 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1364 are shorted:
* D1364 12 12 D_lateral AREA=2.3749375f    ; (-1733.5 -1166 -1699.5 -1162)CMOSN1364 12 12 D_lateral AREA=2.3749375f    
C1357 386 12  184.041f    ; (1836.5 -1227 2122.5 -941)CMOSN.041f    
M1356 644 642 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M1355 644 642 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D1354 are shorted:
* D1354 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1218 1670.5 -1214)CMOSN1354 12 12 D_lateral AREA=2.5E-016    
M1353 644 642 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M1352 644 642 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
* Pins of element D1351 are shorted:
* D1351 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1218 1542.5 -1214)CMOSN1351 8 8 D_lateral AREA=2.5E-016    
M1350 442 683 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M1349 8 683 442 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
* Pins of element D1348 are shorted:
* D1348 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1214 -1605.499 -1210)CMOSN1348 8 8 D_lateral AREA=2.5E-016    
M1347 442 683 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M1346 442 683 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D1345 are shorted:
* D1345 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1214 -1733.499 -1210)CMOSN1345 12 12 D_lateral AREA=2.5E-016    
C1342 684 12  184.041f    ; (-2185.5 -1223 -1899.5 -937)CMOSN.041f    
M1333 685 690 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1332 685 690 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D1331 are shorted:
* D1331 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1404 1697.5 -1400)CMOSN1331 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1330 are shorted:
* D1330 12 12 D_lateral AREA=3.249875f    ; (1661.5 -1388 1697.5 -1380)CMOSN1330 12 12 D_lateral AREA=3.249875f    
* Pins of element D1329 are shorted:
* D1329 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1401 1637.501 -1397)CMOSN1329 8 8 D_lateral AREA=2.5E-016    
M1327 685 686 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1325 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1323 685 686 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1320 685 686 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1319 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1318 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D1317 are shorted:
* D1317 8 8 D_lateral AREA=8.875125f    ; (1502.499 -1385 1637.501 -1380.999)CMOSN1317 8 8 D_lateral AREA=8.875125f    
M1312 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1310 8 689 688 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1308 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1305 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1304 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1303 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1302 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1301 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1300 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D1299 are shorted:
* D1299 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1400 -1760.499 -1396)CMOSN1299 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1298 are shorted:
* D1298 12 12 D_lateral AREA=3.249875f    ; (-1760.5 -1384 -1724.5 -1376)CMOSN1298 12 12 D_lateral AREA=3.249875f    
* Pins of element D1297 are shorted:
* D1297 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -1397 -1700.5 -1393)CMOSN1297 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1296 are shorted:
* D1296 8 8 D_lateral AREA=8.875125f    ; (-1700.501 -1381 -1565.499 -1376.999)CMOSN1296 8 8 D_lateral AREA=8.875125f    
M1283 686 8 690 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M1282 690 8 686 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M1281 686 8 690 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M1280 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1279 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1278 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1277 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1276 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1275 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1274 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1273 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1272 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1271 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1270 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1269 12 690 685 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M1268 685 690 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D1267 are shorted:
* D1267 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1500 1697.5 -1496)CMOSN1267 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1266 are shorted:
* D1266 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1484 1697.5 -1480)CMOSN1266 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1265 are shorted:
* D1265 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1468 1697.5 -1464)CMOSN1265 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1264 are shorted:
* D1264 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1452 1697.5 -1448)CMOSN1264 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1263 are shorted:
* D1263 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1436 1697.5 -1432)CMOSN1263 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1262 are shorted:
* D1262 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1420 1697.5 -1416)CMOSN1262 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1261 are shorted:
* D1261 8 8 D_lateral AREA=1.8125625f    ; (1614.5 -1451.001 1637.501 -1445)CMOSN1261 8 8 D_lateral AREA=1.8125625f    
* Pins of element D1260 are shorted:
* D1260 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1433 1637.501 -1429)CMOSN1260 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1259 are shorted:
* D1259 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1417 1637.501 -1413)CMOSN1259 8 8 D_lateral AREA=2.5E-016    
M1257 686 403 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M1256 686 403 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M1255 686 403 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M1254 686 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M1253 8 686 685 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1251 685 686 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1249 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1247 685 686 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1245 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D1242 are shorted:
* D1242 8 8 D_lateral AREA=2.5E-016    ; (1558.499 -1492 1558.5 -1488)CMOSN1242 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1241 are shorted:
* D1241 8 8 D_lateral AREA=3.5625625f    ; (1558.499 -1476 1605.5 -1465.999)CMOSN1241 8 8 D_lateral AREA=3.5625625f    
M1240 8 686 685 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1239 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1238 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1237 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1236 8 686 685 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1230 8 12 689 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M1229 689 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M1228 689 12 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M1227 689 12 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
M1226 8 689 688 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1224 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1222 8 689 688 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1220 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1218 8 689 688 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D1215 are shorted:
* D1215 8 8 D_lateral AREA=2.5E-016    ; (-1621.5 -1488 -1621.499 -1484)CMOSN1215 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1214 are shorted:
* D1214 8 8 D_lateral AREA=3.5625625f    ; (-1668.5 -1472 -1621.499 -1461.999)CMOSN1214 8 8 D_lateral AREA=3.5625625f    
* Pins of element D1213 are shorted:
* D1213 8 8 D_lateral AREA=3.125E-016    ; (-1621.5 -1505 -1621.499 -1500)CMOSN1213 8 8 D_lateral AREA=3.125E-016    
* Pins of element D1212 are shorted:
* D1212 8 8 D_lateral AREA=3.125E-016    ; (-1674.501 -1505 -1674.5 -1500)CMOSN1212 8 8 D_lateral AREA=3.125E-016    
M1211 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M1210 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1209 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1208 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1207 688 689 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1206 693 12 689 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M1205 689 12 693 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M1204 693 12 689 12 CMOSN L=500n W=3.25u AD=2.53125p PD=5u AS=4.875p PS=9.5u    
M1202 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1201 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1200 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1199 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1198 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1197 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1196 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1195 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1194 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1193 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1192 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1191 688 693 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D1190 are shorted:
* D1190 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1496 -1760.499 -1492)CMOSN1190 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1189 are shorted:
* D1189 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1480 -1760.499 -1476)CMOSN1189 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1188 are shorted:
* D1188 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1464 -1760.499 -1460)CMOSN1188 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1187 are shorted:
* D1187 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1448 -1760.499 -1444)CMOSN1187 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1186 are shorted:
* D1186 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1432 -1760.499 -1428)CMOSN1186 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1185 are shorted:
* D1185 12 12 D_lateral AREA=2.5E-016    ; (-1760.5 -1416 -1760.499 -1412)CMOSN1185 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1184 are shorted:
* D1184 8 8 D_lateral AREA=1.8125625f    ; (-1700.501 -1447.001 -1677.5 -1441)CMOSN1184 8 8 D_lateral AREA=1.8125625f    
* Pins of element D1183 are shorted:
* D1183 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -1429 -1700.5 -1425)CMOSN1183 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1182 are shorted:
* D1182 8 8 D_lateral AREA=2.5E-016    ; (-1700.501 -1413 -1700.5 -1409)CMOSN1182 8 8 D_lateral AREA=2.5E-016    
M1174 685 690 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1173 690 403 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1172 12 403 690 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1171 690 403 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M1170 690 691 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M1169 691 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M1168 692 685 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M1167 692 685 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D1166 are shorted:
* D1166 12 12 D_lateral AREA=2f    ; (1641.499 -1551 1651.5 -1539)CMOSN1166 12 12 D_lateral AREA=2f    
* Pins of element D1165 are shorted:
* D1165 12 12 D_lateral AREA=2.687375f    ; (1634.5 -1598 1669.5 -1594)CMOSN1165 12 12 D_lateral AREA=2.687375f    
* Pins of element D1164 are shorted:
* D1164 12 12 D_lateral AREA=2.4374375f    ; (1634.5 -1582 1667.5 -1576)CMOSN1164 12 12 D_lateral AREA=2.4374375f    
* Pins of element D1163 are shorted:
* D1163 12 12 D_lateral AREA=2.3749375f    ; (1663.5 -1516 1697.5 -1512)CMOSN1163 12 12 D_lateral AREA=2.3749375f    
* Pins of element D1161 are shorted:
* D1161 12 12 D_lateral AREA=3.75E-016    ; (1632.5 -1548 1632.501 -1542)CMOSN1161 12 12 D_lateral AREA=3.75E-016    
* Pins of element D1159 are shorted:
* D1159 8 8 D_lateral AREA=3.125E-016    ; (1611.5 -1509 1611.501 -1504)CMOSN1159 8 8 D_lateral AREA=3.125E-016    
M1158 692 685 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1157 692 685 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M1156 690 691 686 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M1155 686 691 690 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M1154 690 691 686 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M1153 691 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D1152 are shorted:
* D1152 8 8 D_lateral AREA=4.1250625f    ; (1552.5 -1582 1610.501 -1573.999)CMOSN1152 8 8 D_lateral AREA=4.1250625f    
* Pins of element D1151 are shorted:
* D1151 8 8 D_lateral AREA=4.375E-016    ; (1610.5 -1602 1610.501 -1595)CMOSN1151 8 8 D_lateral AREA=4.375E-016    
* Pins of element D1149 are shorted:
* D1149 8 8 D_lateral AREA=4.062625f    ; (1558.499 -1564.001 1611.501 -1558)CMOSN1149 8 8 D_lateral AREA=4.062625f    
* Pins of element D1148 are shorted:
* D1148 8 8 D_lateral AREA=3.125E-016    ; (1558.499 -1509 1558.5 -1504)CMOSN1148 8 8 D_lateral AREA=3.125E-016    
M1147 696 697 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1146 697 688 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M1145 697 688 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
M1144 693 694 689 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M1143 689 694 693 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M1142 693 694 689 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M1141 694 12 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D1140 are shorted:
* D1140 8 8 D_lateral AREA=8.625f    ; (-1668.5 -1602 -1605.499 -1590)CMOSN1140 8 8 D_lateral AREA=8.625f    
* Pins of element D1139 are shorted:
* D1139 8 8 D_lateral AREA=4.375E-016    ; (-1673.501 -1598 -1673.5 -1591)CMOSN1139 8 8 D_lateral AREA=4.375E-016    
* Pins of element D1138 are shorted:
* D1138 8 8 D_lateral AREA=4.1250625f    ; (-1673.501 -1578 -1615.5 -1569.999)CMOSN1138 8 8 D_lateral AREA=4.1250625f    
* Pins of element D1137 are shorted:
* D1137 8 8 D_lateral AREA=4.062625f    ; (-1674.501 -1560.001 -1621.499 -1554)CMOSN1137 8 8 D_lateral AREA=4.062625f    
M1136 12 693 688 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M1135 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M1134 693 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1133 12 12 693 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M1132 693 12 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M1131 693 694 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M1130 694 12 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M1129 697 688 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M1128 697 688 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D1127 are shorted:
* D1127 12 12 D_lateral AREA=3.75E-016    ; (-1695.501 -1544 -1695.5 -1538)CMOSN1127 12 12 D_lateral AREA=3.75E-016    
* Pins of element D1126 are shorted:
* D1126 12 12 D_lateral AREA=2f    ; (-1714.5 -1547 -1704.499 -1535)CMOSN1126 12 12 D_lateral AREA=2f    
* Pins of element D1125 are shorted:
* D1125 12 12 D_lateral AREA=2.4374375f    ; (-1730.5 -1578 -1697.5 -1572)CMOSN1125 12 12 D_lateral AREA=2.4374375f    
* Pins of element D1124 are shorted:
* D1124 12 12 D_lateral AREA=2.687375f    ; (-1732.5 -1594 -1697.5 -1590)CMOSN1124 12 12 D_lateral AREA=2.687375f    
* Pins of element D1123 are shorted:
* D1123 12 12 D_lateral AREA=2.3749375f    ; (-1760.5 -1512 -1726.5 -1508)CMOSN1123 12 12 D_lateral AREA=2.3749375f    
* Pins of element D1122 are shorted:
* D1122 12 12 D_lateral AREA=2.3749375f    ; (-1733.5 -1602 -1699.5 -1598)CMOSN1122 12 12 D_lateral AREA=2.3749375f    
C1115 685 12  184.041f    ; (1836.5 -1663 2122.5 -1377)CMOSN.041f    
M1114 695 692 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M1113 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1112 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1111 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1110 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1109 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1108 695 692 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
* Pins of element D1107 are shorted:
* D1107 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1654 1670.5 -1650)CMOSN1107 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1106 are shorted:
* D1106 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1638 1670.5 -1634)CMOSN1106 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1105 are shorted:
* D1105 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -1622 1670.5 -1618)CMOSN1105 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1104 are shorted:
* D1104 12 12 D_lateral AREA=2.3749375f    ; (1636.5 -1606 1670.5 -1602)CMOSN1104 12 12 D_lateral AREA=2.3749375f    
M1103 695 692 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M1102 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1101 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1100 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1099 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1098 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1097 695 692 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
* Pins of element D1096 are shorted:
* D1096 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1654 1542.5 -1650)CMOSN1096 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1095 are shorted:
* D1095 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1638 1542.5 -1634)CMOSN1095 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1094 are shorted:
* D1094 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -1622 1542.5 -1618)CMOSN1094 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1093 are shorted:
* D1093 8 8 D_lateral AREA=8.625f    ; (1542.499 -1606 1605.5 -1594)CMOSN1093 8 8 D_lateral AREA=8.625f    
M1092 696 697 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M1091 8 697 696 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M1090 696 697 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1089 8 697 696 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M1088 696 697 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M1087 8 697 696 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
* Pins of element D1086 are shorted:
* D1086 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1650 -1605.499 -1646)CMOSN1086 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1085 are shorted:
* D1085 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1634 -1605.499 -1630)CMOSN1085 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1084 are shorted:
* D1084 8 8 D_lateral AREA=2.5E-016    ; (-1605.5 -1618 -1605.499 -1614)CMOSN1084 8 8 D_lateral AREA=2.5E-016    
M1083 696 697 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M1082 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1081 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1080 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1079 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1078 696 697 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D1077 are shorted:
* D1077 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1650 -1733.499 -1646)CMOSN1077 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1076 are shorted:
* D1076 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1634 -1733.499 -1630)CMOSN1076 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1075 are shorted:
* D1075 12 12 D_lateral AREA=2.5E-016    ; (-1733.5 -1618 -1733.499 -1614)CMOSN1075 12 12 D_lateral AREA=2.5E-016    
C1072 688 12  184.041f    ; (-2185.5 -1659 -1899.5 -1373)CMOSN.041f    
M1058 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1057 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1056 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1055 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1054 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1053 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1052 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1051 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1050 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M1049 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
* Pins of element D1048 are shorted:
* D1048 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1904 1697.5 -1900)CMOSN1048 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1047 are shorted:
* D1047 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1888 1697.5 -1884)CMOSN1047 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1046 are shorted:
* D1046 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1872 1697.5 -1868)CMOSN1046 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1045 are shorted:
* D1045 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1856 1697.5 -1852)CMOSN1045 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1044 are shorted:
* D1044 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1840 1697.5 -1836)CMOSN1044 12 12 D_lateral AREA=2.5E-016    
* Pins of element D1043 are shorted:
* D1043 12 12 D_lateral AREA=3.249875f    ; (1661.5 -1824 1697.5 -1816)CMOSN1043 12 12 D_lateral AREA=3.249875f    
* Pins of element D1042 are shorted:
* D1042 8 8 D_lateral AREA=1.8125625f    ; (1614.5 -1887.001 1637.501 -1881)CMOSN1042 8 8 D_lateral AREA=1.8125625f    
* Pins of element D1041 are shorted:
* D1041 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1869 1637.501 -1865)CMOSN1041 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1040 are shorted:
* D1040 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1853 1637.501 -1849)CMOSN1040 8 8 D_lateral AREA=2.5E-016    
* Pins of element D1039 are shorted:
* D1039 8 8 D_lateral AREA=2.5E-016    ; (1637.5 -1837 1637.501 -1833)CMOSN1039 8 8 D_lateral AREA=2.5E-016    
M1037 8 701 700 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1035 700 701 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1033 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1031 700 701 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1029 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1027 700 701 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M1025 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1023 700 701 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1019 700 701 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M1018 8 701 700 8 CMOSP L=500n W=16u AD=25p PD=35.5u AS=12p PS=17.5u    
M1017 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1016 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1015 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1014 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1013 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M1012 8 701 700 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
* Pins of element D1011 are shorted:
* D1011 8 8 D_lateral AREA=8.875125f    ; (1502.499 -1821 1637.501 -1816.999)CMOSN1011 8 8 D_lateral AREA=8.875125f    
M1003 701 8 702 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M1002 702 8 701 12 CMOSN L=500n W=3.5u AD=5.25p PD=10u AS=2.625p PS=5u    
M1001 701 8 702 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=2.53125p PS=5u    
M1000 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M999 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M998 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M997 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M996 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M995 700 702 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M994 702 537 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M993 12 537 702 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M992 702 537 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M991 702 703 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M990 703 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
* Pins of element D989 are shorted:
* D989 12 12 D_lateral AREA=2f    ; (1641.499 -1987 1651.5 -1975)CMOSN989 12 12 D_lateral AREA=2f    
* Pins of element D988 are shorted:
* D988 12 12 D_lateral AREA=2.3749375f    ; (1663.5 -1952 1697.5 -1948)CMOSN988 12 12 D_lateral AREA=2.3749375f    
* Pins of element D987 are shorted:
* D987 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1936 1697.5 -1932)CMOSN987 12 12 D_lateral AREA=2.5E-016    
* Pins of element D986 are shorted:
* D986 12 12 D_lateral AREA=2.5E-016    ; (1697.499 -1920 1697.5 -1916)CMOSN986 12 12 D_lateral AREA=2.5E-016    
* Pins of element D985 are shorted:
* D985 12 12 D_lateral AREA=3.75E-016    ; (1632.5 -1984 1632.501 -1978)CMOSN985 12 12 D_lateral AREA=3.75E-016    
* Pins of element D983 are shorted:
* D983 8 8 D_lateral AREA=3.125E-016    ; (1611.5 -1945 1611.501 -1940)CMOSN983 8 8 D_lateral AREA=3.125E-016    
M982 701 537 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M981 701 537 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=9.0625p PS=14u    
M980 701 537 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M979 702 703 701 8 CMOSP L=500n W=11.75u AD=17.125p PD=26.5u AS=8.8125p PS=13.25u    
M978 701 703 702 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M977 702 703 701 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.625p PS=26.5u    
M976 703 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M975 701 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
* Pins of element D974 are shorted:
* D974 8 8 D_lateral AREA=4.062625f    ; (1558.499 -2000.001 1611.501 -1994)CMOSN974 8 8 D_lateral AREA=4.062625f    
* Pins of element D973 are shorted:
* D973 8 8 D_lateral AREA=3.125E-016    ; (1558.499 -1945 1558.5 -1940)CMOSN973 8 8 D_lateral AREA=3.125E-016    
* Pins of element D972 are shorted:
* D972 8 8 D_lateral AREA=2.5E-016    ; (1558.499 -1928 1558.5 -1924)CMOSN972 8 8 D_lateral AREA=2.5E-016    
* Pins of element D971 are shorted:
* D971 8 8 D_lateral AREA=3.5625625f    ; (1558.499 -1912 1605.5 -1901.999)CMOSN971 8 8 D_lateral AREA=3.5625625f    
C964 700 12  184.041f    ; (1836.5 -2099 2122.5 -1813)CMOSN.041f    
M963 705 704 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
M962 12 704 705 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M961 705 704 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M960 12 704 705 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M959 705 704 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M958 12 704 705 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M957 705 704 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M956 704 700 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
M955 704 700 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D954 are shorted:
* D954 12 12 D_lateral AREA=2.687375f    ; (1634.5 -2034 1669.5 -2030)CMOSN954 12 12 D_lateral AREA=2.687375f    
* Pins of element D953 are shorted:
* D953 12 12 D_lateral AREA=2.4374375f    ; (1634.5 -2018 1667.5 -2012)CMOSN953 12 12 D_lateral AREA=2.4374375f    
* Pins of element D952 are shorted:
* D952 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -2090 1670.5 -2086)CMOSN952 12 12 D_lateral AREA=2.5E-016    
* Pins of element D951 are shorted:
* D951 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -2074 1670.5 -2070)CMOSN951 12 12 D_lateral AREA=2.5E-016    
* Pins of element D950 are shorted:
* D950 12 12 D_lateral AREA=2.5E-016    ; (1670.499 -2058 1670.5 -2054)CMOSN950 12 12 D_lateral AREA=2.5E-016    
* Pins of element D949 are shorted:
* D949 12 12 D_lateral AREA=2.3749375f    ; (1636.5 -2042 1670.5 -2038)CMOSN949 12 12 D_lateral AREA=2.3749375f    
M948 705 704 8 8 CMOSP L=500n W=16u AD=24p PD=35u AS=12.25p PS=18u    
M947 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M946 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M945 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M944 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M943 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M942 705 704 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M941 704 700 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M940 704 700 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=35.5p PS=37.5u    
* Pins of element D939 are shorted:
* D939 8 8 D_lateral AREA=4.1250625f    ; (1552.5 -2018 1610.501 -2009.999)CMOSN939 8 8 D_lateral AREA=4.1250625f    
* Pins of element D938 are shorted:
* D938 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -2090 1542.5 -2086)CMOSN938 8 8 D_lateral AREA=2.5E-016    
* Pins of element D937 are shorted:
* D937 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -2074 1542.5 -2070)CMOSN937 8 8 D_lateral AREA=2.5E-016    
* Pins of element D936 are shorted:
* D936 8 8 D_lateral AREA=2.5E-016    ; (1542.499 -2058 1542.5 -2054)CMOSN936 8 8 D_lateral AREA=2.5E-016    
* Pins of element D935 are shorted:
* D935 8 8 D_lateral AREA=4.375E-016    ; (1610.5 -2038 1610.501 -2031)CMOSN935 8 8 D_lateral AREA=4.375E-016    
* Pins of element D934 are shorted:
* D934 8 8 D_lateral AREA=8.625f    ; (1542.499 -2042 1605.5 -2030)CMOSN934 8 8 D_lateral AREA=8.625f    
C931 8 12  184.041f    ; (-2185.5 -2095 -1899.5 -1809)CMOSN.041f    
M865 8 8 714 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M863 8 714 706 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M861 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M859 8 714 706 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M857 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M855 8 714 706 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M853 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M851 8 714 706 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M849 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D847 are shorted:
* D847 8 8 D_lateral AREA=3.5625625f    ; (1320.5 -2285 1330.501 -2237.999)CMOSN847 8 8 D_lateral AREA=3.5625625f    
M846 8 536 714 8 CMOSP L=500n W=11.5u AD=9.0625p PD=14u AS=8.90625p PS=13.75u    
M845 8 536 714 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M844 714 536 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M843 8 706 717 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M842 714 715 716 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M841 716 715 714 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M840 714 715 716 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M839 715 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D838 are shorted:
* D838 8 8 D_lateral AREA=4.1250625f    ; (1214.5 -2290.001 1222.501 -2232)CMOSN838 8 8 D_lateral AREA=4.1250625f    
* Pins of element D837 are shorted:
* D837 8 8 D_lateral AREA=2.5E-016    ; (1304.5 -2238 1308.5 -2237.999)CMOSN837 8 8 D_lateral AREA=2.5E-016    
* Pins of element D836 are shorted:
* D836 8 8 D_lateral AREA=3.125E-016    ; (1287.5 -2291.001 1292.5 -2291)CMOSN836 8 8 D_lateral AREA=3.125E-016    
* Pins of element D835 are shorted:
* D835 8 8 D_lateral AREA=3.125E-016    ; (1287.5 -2238 1292.5 -2237.999)CMOSN835 8 8 D_lateral AREA=3.125E-016    
* Pins of element D834 are shorted:
* D834 8 8 D_lateral AREA=4.062625f    ; (1232.499 -2291.001 1238.5 -2237.999)CMOSN834 8 8 D_lateral AREA=4.062625f    
M833 8 717 718 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M832 718 717 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M831 8 717 718 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M830 718 717 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M829 8 717 718 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M828 718 717 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M827 8 717 718 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M826 717 706 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
* Pins of element D825 are shorted:
* D825 8 8 D_lateral AREA=4.375E-016    ; (1194.5 -2290.001 1201.5 -2290)CMOSN825 8 8 D_lateral AREA=4.375E-016    
* Pins of element D824 are shorted:
* D824 8 8 D_lateral AREA=8.625f    ; (1190.5 -2285 1202.5 -2221.999)CMOSN824 8 8 D_lateral AREA=8.625f    
* Pins of element D823 are shorted:
* D823 8 8 D_lateral AREA=2.5E-016    ; (1174.5 -2222 1178.5 -2221.999)CMOSN823 8 8 D_lateral AREA=2.5E-016    
* Pins of element D822 are shorted:
* D822 8 8 D_lateral AREA=2.5E-016    ; (1158.5 -2222 1162.5 -2221.999)CMOSN822 8 8 D_lateral AREA=2.5E-016    
* Pins of element D821 are shorted:
* D821 8 8 D_lateral AREA=2.5E-016    ; (1142.5 -2222 1146.5 -2221.999)CMOSN821 8 8 D_lateral AREA=2.5E-016    
M819 8 720 723 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M817 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M815 8 720 723 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M813 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M811 8 720 723 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M809 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M807 8 720 723 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M805 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M803 720 698 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M802 8 698 720 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M801 720 698 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M800 720 721 719 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M799 719 721 720 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M798 720 721 719 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M797 8 8 720 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
* Pins of element D795 are shorted:
* D795 8 8 D_lateral AREA=3.5625625f    ; (884.5 -2285 894.501 -2237.999)CMOSN795 8 8 D_lateral AREA=3.5625625f    
* Pins of element D794 are shorted:
* D794 8 8 D_lateral AREA=2.5E-016    ; (868.5 -2238 872.5 -2237.999)CMOSN794 8 8 D_lateral AREA=2.5E-016    
* Pins of element D793 are shorted:
* D793 8 8 D_lateral AREA=3.125E-016    ; (851.5 -2291.001 856.5 -2291)CMOSN793 8 8 D_lateral AREA=3.125E-016    
* Pins of element D792 are shorted:
* D792 8 8 D_lateral AREA=3.125E-016    ; (851.5 -2238 856.5 -2237.999)CMOSN792 8 8 D_lateral AREA=3.125E-016    
M791 8 707 722 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M790 722 707 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M789 8 707 722 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M788 722 707 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M787 8 707 722 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M786 722 707 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M785 8 723 707 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M784 707 723 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M783 721 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D782 are shorted:
* D782 8 8 D_lateral AREA=4.1250625f    ; (778.5 -2290.001 786.501 -2232)CMOSN782 8 8 D_lateral AREA=4.1250625f    
* Pins of element D781 are shorted:
* D781 8 8 D_lateral AREA=4.375E-016    ; (758.5 -2290.001 765.5 -2290)CMOSN781 8 8 D_lateral AREA=4.375E-016    
* Pins of element D780 are shorted:
* D780 8 8 D_lateral AREA=8.625f    ; (754.5 -2285 766.5 -2221.999)CMOSN780 8 8 D_lateral AREA=8.625f    
* Pins of element D779 are shorted:
* D779 8 8 D_lateral AREA=2.5E-016    ; (738.5 -2222 742.5 -2221.999)CMOSN779 8 8 D_lateral AREA=2.5E-016    
* Pins of element D778 are shorted:
* D778 8 8 D_lateral AREA=2.5E-016    ; (722.5 -2222 726.5 -2221.999)CMOSN778 8 8 D_lateral AREA=2.5E-016    
* Pins of element D777 are shorted:
* D777 8 8 D_lateral AREA=4.062625f    ; (796.499 -2291.001 802.5 -2237.999)CMOSN777 8 8 D_lateral AREA=4.062625f    
M776 8 707 722 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
* Pins of element D775 are shorted:
* D775 8 8 D_lateral AREA=2.5E-016    ; (706.5 -2222 710.5 -2221.999)CMOSN775 8 8 D_lateral AREA=2.5E-016    
M773 8 724 727 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M771 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M769 8 724 727 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M767 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M765 724 699 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M764 8 699 724 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M763 724 699 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M762 8 8 724 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M760 8 724 727 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M758 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M756 8 724 727 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M754 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D752 are shorted:
* D752 8 8 D_lateral AREA=3.5625625f    ; (448.5 -2285 458.501 -2237.999)CMOSN752 8 8 D_lateral AREA=3.5625625f    
* Pins of element D751 are shorted:
* D751 8 8 D_lateral AREA=2.5E-016    ; (432.5 -2238 436.5 -2237.999)CMOSN751 8 8 D_lateral AREA=2.5E-016    
* Pins of element D750 are shorted:
* D750 8 8 D_lateral AREA=3.125E-016    ; (415.5 -2291.001 420.5 -2291)CMOSN750 8 8 D_lateral AREA=3.125E-016    
* Pins of element D749 are shorted:
* D749 8 8 D_lateral AREA=3.125E-016    ; (415.5 -2238 420.5 -2237.999)CMOSN749 8 8 D_lateral AREA=3.125E-016    
M748 8 709 708 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M747 8 727 709 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M746 709 727 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M745 724 726 725 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M744 725 726 724 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M743 724 726 725 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M742 726 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D741 are shorted:
* D741 8 8 D_lateral AREA=4.1250625f    ; (342.5 -2290.001 350.501 -2232)CMOSN741 8 8 D_lateral AREA=4.1250625f    
* Pins of element D740 are shorted:
* D740 8 8 D_lateral AREA=4.375E-016    ; (322.5 -2290.001 329.5 -2290)CMOSN740 8 8 D_lateral AREA=4.375E-016    
* Pins of element D739 are shorted:
* D739 8 8 D_lateral AREA=8.625f    ; (318.5 -2285 330.5 -2221.999)CMOSN739 8 8 D_lateral AREA=8.625f    
* Pins of element D738 are shorted:
* D738 8 8 D_lateral AREA=4.062625f    ; (360.499 -2291.001 366.5 -2237.999)CMOSN738 8 8 D_lateral AREA=4.062625f    
M737 708 709 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M736 8 709 708 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M735 708 709 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M734 8 709 708 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M733 708 709 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M732 8 709 708 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
* Pins of element D731 are shorted:
* D731 8 8 D_lateral AREA=2.5E-016    ; (302.5 -2222 306.5 -2221.999)CMOSN731 8 8 D_lateral AREA=2.5E-016    
* Pins of element D730 are shorted:
* D730 8 8 D_lateral AREA=2.5E-016    ; (286.5 -2222 290.5 -2221.999)CMOSN730 8 8 D_lateral AREA=2.5E-016    
* Pins of element D729 are shorted:
* D729 8 8 D_lateral AREA=2.5E-016    ; (270.5 -2222 274.5 -2221.999)CMOSN729 8 8 D_lateral AREA=2.5E-016    
M726 8 728 710 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M724 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M722 8 728 710 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M720 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M718 8 728 710 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M716 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M714 8 728 710 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M712 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D709 are shorted:
* D709 8 8 D_lateral AREA=3.5625625f    ; (12.5 -2285 22.501 -2237.999)CMOSN709 8 8 D_lateral AREA=3.5625625f    
M708 728 687 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M707 8 687 728 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M706 728 687 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M705 728 730 729 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M704 729 730 728 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M703 728 730 729 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M702 730 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M701 728 8 8 8 CMOSP L=500n W=12.25u AD=8.90625p PD=13.75u AS=33.4375p PS=31u    
* Pins of element D699 are shorted:
* D699 8 8 D_lateral AREA=2.5E-016    ; (-3.5 -2238 0.5 -2237.999)CMOSN699 8 8 D_lateral AREA=2.5E-016    
* Pins of element D698 are shorted:
* D698 8 8 D_lateral AREA=3.125E-016    ; (-20.5 -2291.001 -15.5 -2291)CMOSN698 8 8 D_lateral AREA=3.125E-016    
* Pins of element D697 are shorted:
* D697 8 8 D_lateral AREA=3.125E-016    ; (-20.5 -2238 -15.5 -2237.999)CMOSN697 8 8 D_lateral AREA=3.125E-016    
* Pins of element D696 are shorted:
* D696 8 8 D_lateral AREA=4.062625f    ; (-75.501 -2291.001 -69.5 -2237.999)CMOSN696 8 8 D_lateral AREA=4.062625f    
M695 8 731 732 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M694 732 731 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M693 8 731 732 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M692 732 731 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M691 8 731 732 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M690 732 731 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M689 8 731 732 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M688 8 710 731 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M687 731 710 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
* Pins of element D686 are shorted:
* D686 8 8 D_lateral AREA=4.1250625f    ; (-93.5 -2290.001 -85.499 -2232)CMOSN686 8 8 D_lateral AREA=4.1250625f    
* Pins of element D685 are shorted:
* D685 8 8 D_lateral AREA=4.375E-016    ; (-113.5 -2290.001 -106.5 -2290)CMOSN685 8 8 D_lateral AREA=4.375E-016    
* Pins of element D684 are shorted:
* D684 8 8 D_lateral AREA=8.625f    ; (-117.5 -2285 -105.5 -2221.999)CMOSN684 8 8 D_lateral AREA=8.625f    
* Pins of element D683 are shorted:
* D683 8 8 D_lateral AREA=2.5E-016    ; (-133.5 -2222 -129.5 -2221.999)CMOSN683 8 8 D_lateral AREA=2.5E-016    
* Pins of element D682 are shorted:
* D682 8 8 D_lateral AREA=2.5E-016    ; (-149.5 -2222 -145.5 -2221.999)CMOSN682 8 8 D_lateral AREA=2.5E-016    
* Pins of element D681 are shorted:
* D681 8 8 D_lateral AREA=2.5E-016    ; (-165.5 -2222 -161.5 -2221.999)CMOSN681 8 8 D_lateral AREA=2.5E-016    
M679 8 733 711 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M677 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M675 8 733 711 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M673 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M671 8 733 711 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M669 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M667 8 733 711 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M665 733 734 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M664 8 734 733 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M663 733 734 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M662 733 735 712 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M661 712 735 733 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M660 733 735 712 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M659 8 8 733 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M657 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D655 are shorted:
* D655 8 8 D_lateral AREA=3.5625625f    ; (-423.5 -2285 -413.499 -2237.999)CMOSN655 8 8 D_lateral AREA=3.5625625f    
* Pins of element D654 are shorted:
* D654 8 8 D_lateral AREA=2.5E-016    ; (-439.5 -2238 -435.5 -2237.999)CMOSN654 8 8 D_lateral AREA=2.5E-016    
* Pins of element D653 are shorted:
* D653 8 8 D_lateral AREA=3.125E-016    ; (-456.5 -2291.001 -451.5 -2291)CMOSN653 8 8 D_lateral AREA=3.125E-016    
* Pins of element D652 are shorted:
* D652 8 8 D_lateral AREA=3.125E-016    ; (-456.5 -2238 -451.5 -2237.999)CMOSN652 8 8 D_lateral AREA=3.125E-016    
M651 8 713 736 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M650 736 713 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M649 8 713 736 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M648 736 713 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M647 8 713 736 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M646 8 711 713 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M645 713 711 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M644 735 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D643 are shorted:
* D643 8 8 D_lateral AREA=4.1250625f    ; (-529.5 -2290.001 -521.499 -2232)CMOSN643 8 8 D_lateral AREA=4.1250625f    
* Pins of element D642 are shorted:
* D642 8 8 D_lateral AREA=4.375E-016    ; (-549.5 -2290.001 -542.5 -2290)CMOSN642 8 8 D_lateral AREA=4.375E-016    
* Pins of element D641 are shorted:
* D641 8 8 D_lateral AREA=8.625f    ; (-553.5 -2285 -541.5 -2221.999)CMOSN641 8 8 D_lateral AREA=8.625f    
* Pins of element D640 are shorted:
* D640 8 8 D_lateral AREA=2.5E-016    ; (-569.5 -2222 -565.5 -2221.999)CMOSN640 8 8 D_lateral AREA=2.5E-016    
* Pins of element D639 are shorted:
* D639 8 8 D_lateral AREA=2.5E-016    ; (-585.5 -2222 -581.5 -2221.999)CMOSN639 8 8 D_lateral AREA=2.5E-016    
* Pins of element D638 are shorted:
* D638 8 8 D_lateral AREA=4.062625f    ; (-511.501 -2291.001 -505.5 -2237.999)CMOSN638 8 8 D_lateral AREA=4.062625f    
M637 736 713 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M636 8 713 736 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
* Pins of element D635 are shorted:
* D635 8 8 D_lateral AREA=2.5E-016    ; (-601.5 -2222 -597.5 -2221.999)CMOSN635 8 8 D_lateral AREA=2.5E-016    
M633 8 737 743 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M631 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M629 8 737 743 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M627 737 741 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M626 8 741 737 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M625 737 741 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M624 8 8 737 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
M622 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M620 8 737 743 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M618 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M616 8 737 743 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M614 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
* Pins of element D612 are shorted:
* D612 8 8 D_lateral AREA=3.5625625f    ; (-859.5 -2285 -849.499 -2237.999)CMOSN612 8 8 D_lateral AREA=3.5625625f    
* Pins of element D611 are shorted:
* D611 8 8 D_lateral AREA=2.5E-016    ; (-875.5 -2238 -871.5 -2237.999)CMOSN611 8 8 D_lateral AREA=2.5E-016    
M608 8 743 738 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M607 738 743 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
M606 737 740 739 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M605 739 740 737 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M604 737 740 739 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M603 740 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
* Pins of element D602 are shorted:
* D602 8 8 D_lateral AREA=4.1250625f    ; (-965.5 -2290.001 -957.499 -2232)CMOSN602 8 8 D_lateral AREA=4.1250625f    
* Pins of element D601 are shorted:
* D601 8 8 D_lateral AREA=4.375E-016    ; (-985.5 -2290.001 -978.5 -2290)CMOSN601 8 8 D_lateral AREA=4.375E-016    
* Pins of element D599 are shorted:
* D599 8 8 D_lateral AREA=3.125E-016    ; (-892.5 -2291.001 -887.5 -2291)CMOSN599 8 8 D_lateral AREA=3.125E-016    
* Pins of element D598 are shorted:
* D598 8 8 D_lateral AREA=3.125E-016    ; (-892.5 -2238 -887.5 -2237.999)CMOSN598 8 8 D_lateral AREA=3.125E-016    
* Pins of element D597 are shorted:
* D597 8 8 D_lateral AREA=4.062625f    ; (-947.501 -2291.001 -941.5 -2237.999)CMOSN597 8 8 D_lateral AREA=4.062625f    
M596 8 738 742 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M595 742 738 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M594 8 738 742 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M593 742 738 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M592 8 738 742 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M591 742 738 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M590 8 738 742 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
* Pins of element D589 are shorted:
* D589 8 8 D_lateral AREA=8.625f    ; (-989.5 -2285 -977.5 -2221.999)CMOSN589 8 8 D_lateral AREA=8.625f    
* Pins of element D588 are shorted:
* D588 8 8 D_lateral AREA=2.5E-016    ; (-1005.5 -2222 -1001.5 -2221.999)CMOSN588 8 8 D_lateral AREA=2.5E-016    
* Pins of element D587 are shorted:
* D587 8 8 D_lateral AREA=2.5E-016    ; (-1021.5 -2222 -1017.5 -2221.999)CMOSN587 8 8 D_lateral AREA=2.5E-016    
* Pins of element D586 are shorted:
* D586 8 8 D_lateral AREA=2.5E-016    ; (-1037.5 -2222 -1033.5 -2221.999)CMOSN586 8 8 D_lateral AREA=2.5E-016    
M584 8 744 750 8 CMOSP L=500n W=16u AD=20.8125p PD=35.25u AS=12p PS=17.5u    
M582 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M580 8 744 750 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M578 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M576 8 744 750 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M574 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M572 8 744 750 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M570 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M566 744 747 8 8 CMOSP L=500n W=11.5u AD=8.90625p PD=13.75u AS=9.0625p PS=14u    
M565 8 747 744 8 CMOSP L=500n W=12u AD=9.0625p PD=14u AS=9p PS=13.5u    
M564 744 747 8 8 CMOSP L=500n W=12u AD=9p PD=13.5u AS=19.5625p PS=29.5u    
M563 744 746 745 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=8.8125p PS=13.25u    
M562 745 746 744 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=8.8125p PS=13.25u    
M561 744 746 745 8 CMOSP L=500n W=11.75u AD=8.8125p PD=13.25u AS=17.125p PS=26.5u    
M560 746 8 8 8 CMOSP L=500n W=11.75u AD=17.625p PD=26.5u AS=22.8125p PS=30u    
M559 8 8 744 8 CMOSP L=500n W=12.25u AD=33.4375p PD=31u AS=8.90625p PS=13.75u    
* Pins of element D558 are shorted:
* D558 8 8 D_lateral AREA=3.5625625f    ; (-1295.5 -2285 -1285.499 -2237.999)CMOSN558 8 8 D_lateral AREA=3.5625625f    
* Pins of element D557 are shorted:
* D557 8 8 D_lateral AREA=2.5E-016    ; (-1311.5 -2238 -1307.5 -2237.999)CMOSN557 8 8 D_lateral AREA=2.5E-016    
* Pins of element D556 are shorted:
* D556 8 8 D_lateral AREA=3.125E-016    ; (-1328.5 -2291.001 -1323.5 -2291)CMOSN556 8 8 D_lateral AREA=3.125E-016    
* Pins of element D555 are shorted:
* D555 8 8 D_lateral AREA=3.125E-016    ; (-1328.5 -2238 -1323.5 -2237.999)CMOSN555 8 8 D_lateral AREA=3.125E-016    
* Pins of element D554 are shorted:
* D554 8 8 D_lateral AREA=4.062625f    ; (-1383.501 -2291.001 -1377.5 -2237.999)CMOSN554 8 8 D_lateral AREA=4.062625f    
M553 8 748 749 8 CMOSP L=500n W=16u AD=21.3125p PD=36.25u AS=12p PS=17.5u    
M552 749 748 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M551 8 748 749 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M550 749 748 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M549 8 748 749 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=12p PS=17.5u    
M548 749 748 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.25p PS=18u    
M547 8 748 749 8 CMOSP L=500n W=16u AD=12.25p PD=18u AS=24p PS=35u    
M546 8 750 748 8 CMOSP L=500n W=16u AD=35.5p PD=37.5u AS=12p PS=17.5u    
M545 748 750 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=21.3125p PS=36.25u    
* Pins of element D544 are shorted:
* D544 8 8 D_lateral AREA=4.1250625f    ; (-1401.5 -2290.001 -1393.499 -2232)CMOSN544 8 8 D_lateral AREA=4.1250625f    
* Pins of element D543 are shorted:
* D543 8 8 D_lateral AREA=4.375E-016    ; (-1421.5 -2290.001 -1414.5 -2290)CMOSN543 8 8 D_lateral AREA=4.375E-016    
* Pins of element D542 are shorted:
* D542 8 8 D_lateral AREA=8.625f    ; (-1425.5 -2285 -1413.5 -2221.999)CMOSN542 8 8 D_lateral AREA=8.625f    
* Pins of element D541 are shorted:
* D541 8 8 D_lateral AREA=2.5E-016    ; (-1441.5 -2222 -1437.5 -2221.999)CMOSN541 8 8 D_lateral AREA=2.5E-016    
* Pins of element D540 are shorted:
* D540 8 8 D_lateral AREA=2.5E-016    ; (-1457.5 -2222 -1453.5 -2221.999)CMOSN540 8 8 D_lateral AREA=2.5E-016    
* Pins of element D539 are shorted:
* D539 8 8 D_lateral AREA=2.5E-016    ; (-1473.5 -2222 -1469.5 -2221.999)CMOSN539 8 8 D_lateral AREA=2.5E-016    
* Pins of element D537 are shorted:
* D537 8 8 D_lateral AREA=8.875125f    ; (1411.5 -2317.001 1415.501 -2181.999)CMOSN537 8 8 D_lateral AREA=8.875125f    
M536 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M535 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M534 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M533 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M532 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M531 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M530 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M529 706 714 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M528 714 8 716 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M527 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M526 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M525 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M524 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M523 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M522 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M521 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M520 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M519 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M518 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M517 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M516 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D514 are shorted:
* D514 12 12 D_lateral AREA=3.249875f    ; (1408.5 -2377 1416.5 -2341)CMOSN514 12 12 D_lateral AREA=3.249875f    
* Pins of element D513 are shorted:
* D513 12 12 D_lateral AREA=2.5E-016    ; (1392.5 -2377 1396.5 -2376.999)CMOSN513 12 12 D_lateral AREA=2.5E-016    
* Pins of element D512 are shorted:
* D512 12 12 D_lateral AREA=2.5E-016    ; (1376.5 -2377 1380.5 -2376.999)CMOSN512 12 12 D_lateral AREA=2.5E-016    
* Pins of element D511 are shorted:
* D511 12 12 D_lateral AREA=2.5E-016    ; (1360.5 -2377 1364.5 -2376.999)CMOSN511 12 12 D_lateral AREA=2.5E-016    
* Pins of element D510 are shorted:
* D510 12 12 D_lateral AREA=2.5E-016    ; (1344.5 -2377 1348.5 -2376.999)CMOSN510 12 12 D_lateral AREA=2.5E-016    
* Pins of element D509 are shorted:
* D509 12 12 D_lateral AREA=2.5E-016    ; (1328.5 -2377 1332.5 -2376.999)CMOSN509 12 12 D_lateral AREA=2.5E-016    
* Pins of element D508 are shorted:
* D508 12 12 D_lateral AREA=2.5E-016    ; (1312.5 -2377 1316.5 -2376.999)CMOSN508 12 12 D_lateral AREA=2.5E-016    
* Pins of element D506 are shorted:
* D506 8 8 D_lateral AREA=2.5E-016    ; (1395.5 -2317.001 1399.5 -2317)CMOSN506 8 8 D_lateral AREA=2.5E-016    
* Pins of element D505 are shorted:
* D505 8 8 D_lateral AREA=2.5E-016    ; (1379.5 -2317.001 1383.5 -2317)CMOSN505 8 8 D_lateral AREA=2.5E-016    
* Pins of element D504 are shorted:
* D504 8 8 D_lateral AREA=2.5E-016    ; (1363.5 -2317.001 1367.5 -2317)CMOSN504 8 8 D_lateral AREA=2.5E-016    
* Pins of element D503 are shorted:
* D503 8 8 D_lateral AREA=1.8125625f    ; (1345.499 -2317.001 1351.5 -2294)CMOSN503 8 8 D_lateral AREA=1.8125625f    
M502 716 8 714 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M501 714 8 716 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M500 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M499 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M498 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M497 706 716 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M496 12 536 716 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M495 716 536 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M494 12 536 716 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M493 716 715 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M492 715 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M491 717 706 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
* Pins of element D490 are shorted:
* D490 12 12 D_lateral AREA=3.75E-016    ; (1248.5 -2312.001 1254.5 -2312)CMOSN490 12 12 D_lateral AREA=3.75E-016    
* Pins of element D489 are shorted:
* D489 12 12 D_lateral AREA=2f    ; (1245.5 -2331 1257.5 -2320.999)CMOSN489 12 12 D_lateral AREA=2f    
* Pins of element D488 are shorted:
* D488 12 12 D_lateral AREA=2.4374375f    ; (1214.5 -2347 1220.5 -2314)CMOSN488 12 12 D_lateral AREA=2.4374375f    
* Pins of element D487 are shorted:
* D487 12 12 D_lateral AREA=2.5E-016    ; (1296.5 -2377 1300.5 -2376.999)CMOSN487 12 12 D_lateral AREA=2.5E-016    
* Pins of element D486 are shorted:
* D486 12 12 D_lateral AREA=2.3749375f    ; (1280.5 -2377 1284.5 -2343)CMOSN486 12 12 D_lateral AREA=2.3749375f    
M485 12 717 718 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M484 718 717 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M483 12 717 718 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M482 718 717 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M481 12 717 718 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M480 718 717 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M479 12 717 718 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M478 717 706 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D477 are shorted:
* D477 12 12 D_lateral AREA=2.687375f    ; (1198.5 -2349 1202.5 -2314)CMOSN477 12 12 D_lateral AREA=2.687375f    
* Pins of element D476 are shorted:
* D476 12 12 D_lateral AREA=2.3749375f    ; (1190.5 -2350 1194.5 -2316)CMOSN476 12 12 D_lateral AREA=2.3749375f    
* Pins of element D475 are shorted:
* D475 12 12 D_lateral AREA=2.5E-016    ; (1174.5 -2350 1178.5 -2349.999)CMOSN475 12 12 D_lateral AREA=2.5E-016    
* Pins of element D474 are shorted:
* D474 12 12 D_lateral AREA=2.5E-016    ; (1158.5 -2350 1162.5 -2349.999)CMOSN474 12 12 D_lateral AREA=2.5E-016    
* Pins of element D473 are shorted:
* D473 12 12 D_lateral AREA=2.5E-016    ; (1142.5 -2350 1146.5 -2349.999)CMOSN473 12 12 D_lateral AREA=2.5E-016    
M472 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M471 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M470 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M469 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M468 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M467 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M466 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M465 723 720 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M464 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M463 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M462 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M461 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M460 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M459 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M458 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M457 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D456 are shorted:
* D456 12 12 D_lateral AREA=3.249875f    ; (972.5 -2377 980.5 -2341)CMOSN456 12 12 D_lateral AREA=3.249875f    
* Pins of element D455 are shorted:
* D455 12 12 D_lateral AREA=2.5E-016    ; (956.5 -2377 960.5 -2376.999)CMOSN455 12 12 D_lateral AREA=2.5E-016    
* Pins of element D454 are shorted:
* D454 12 12 D_lateral AREA=2.5E-016    ; (940.5 -2377 944.5 -2376.999)CMOSN454 12 12 D_lateral AREA=2.5E-016    
* Pins of element D453 are shorted:
* D453 12 12 D_lateral AREA=2.5E-016    ; (924.5 -2377 928.5 -2376.999)CMOSN453 12 12 D_lateral AREA=2.5E-016    
* Pins of element D451 are shorted:
* D451 8 8 D_lateral AREA=8.875125f    ; (975.5 -2317.001 979.501 -2181.999)CMOSN451 8 8 D_lateral AREA=8.875125f    
* Pins of element D450 are shorted:
* D450 8 8 D_lateral AREA=2.5E-016    ; (959.5 -2317.001 963.5 -2317)CMOSN450 8 8 D_lateral AREA=2.5E-016    
* Pins of element D449 are shorted:
* D449 8 8 D_lateral AREA=2.5E-016    ; (943.5 -2317.001 947.5 -2317)CMOSN449 8 8 D_lateral AREA=2.5E-016    
* Pins of element D448 are shorted:
* D448 8 8 D_lateral AREA=2.5E-016    ; (927.5 -2317.001 931.5 -2317)CMOSN448 8 8 D_lateral AREA=2.5E-016    
M446 720 8 719 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M445 719 8 720 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M444 720 8 719 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M443 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M442 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M441 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M440 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M439 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M438 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M437 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M436 723 719 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M435 12 698 719 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M434 719 698 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M433 12 698 719 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M432 719 721 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D431 are shorted:
* D431 12 12 D_lateral AREA=3.75E-016    ; (812.5 -2312.001 818.5 -2312)CMOSN431 12 12 D_lateral AREA=3.75E-016    
* Pins of element D429 are shorted:
* D429 12 12 D_lateral AREA=2.5E-016    ; (908.5 -2377 912.5 -2376.999)CMOSN429 12 12 D_lateral AREA=2.5E-016    
* Pins of element D428 are shorted:
* D428 12 12 D_lateral AREA=2.5E-016    ; (892.5 -2377 896.5 -2376.999)CMOSN428 12 12 D_lateral AREA=2.5E-016    
* Pins of element D427 are shorted:
* D427 12 12 D_lateral AREA=2.5E-016    ; (876.5 -2377 880.5 -2376.999)CMOSN427 12 12 D_lateral AREA=2.5E-016    
* Pins of element D426 are shorted:
* D426 12 12 D_lateral AREA=2.5E-016    ; (860.5 -2377 864.5 -2376.999)CMOSN426 12 12 D_lateral AREA=2.5E-016    
* Pins of element D425 are shorted:
* D425 12 12 D_lateral AREA=2.3749375f    ; (844.5 -2377 848.5 -2343)CMOSN425 12 12 D_lateral AREA=2.3749375f    
* Pins of element D424 are shorted:
* D424 8 8 D_lateral AREA=1.8125625f    ; (909.499 -2317.001 915.5 -2294)CMOSN424 8 8 D_lateral AREA=1.8125625f    
M423 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M422 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M421 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M420 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M419 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M418 722 707 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M417 721 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M416 12 723 707 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
M415 707 723 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D414 are shorted:
* D414 12 12 D_lateral AREA=2f    ; (809.5 -2331 821.5 -2320.999)CMOSN414 12 12 D_lateral AREA=2f    
* Pins of element D413 are shorted:
* D413 12 12 D_lateral AREA=2.4374375f    ; (778.5 -2347 784.5 -2314)CMOSN413 12 12 D_lateral AREA=2.4374375f    
* Pins of element D412 are shorted:
* D412 12 12 D_lateral AREA=2.687375f    ; (762.5 -2349 766.5 -2314)CMOSN412 12 12 D_lateral AREA=2.687375f    
* Pins of element D411 are shorted:
* D411 12 12 D_lateral AREA=2.3749375f    ; (754.5 -2350 758.5 -2316)CMOSN411 12 12 D_lateral AREA=2.3749375f    
* Pins of element D410 are shorted:
* D410 12 12 D_lateral AREA=2.5E-016    ; (738.5 -2350 742.5 -2349.999)CMOSN410 12 12 D_lateral AREA=2.5E-016    
* Pins of element D409 are shorted:
* D409 12 12 D_lateral AREA=2.5E-016    ; (722.5 -2350 726.5 -2349.999)CMOSN409 12 12 D_lateral AREA=2.5E-016    
M408 722 707 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
* Pins of element D407 are shorted:
* D407 12 12 D_lateral AREA=2.5E-016    ; (706.5 -2350 710.5 -2349.999)CMOSN407 12 12 D_lateral AREA=2.5E-016    
M406 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M405 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M404 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M403 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M402 727 725 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M401 727 725 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M400 727 725 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D398 are shorted:
* D398 12 12 D_lateral AREA=3.249875f    ; (536.5 -2377 544.5 -2341)CMOSN398 12 12 D_lateral AREA=3.249875f    
* Pins of element D397 are shorted:
* D397 12 12 D_lateral AREA=2.5E-016    ; (520.5 -2377 524.5 -2376.999)CMOSN397 12 12 D_lateral AREA=2.5E-016    
* Pins of element D396 are shorted:
* D396 8 8 D_lateral AREA=8.875125f    ; (539.5 -2317.001 543.501 -2181.999)CMOSN396 8 8 D_lateral AREA=8.875125f    
* Pins of element D395 are shorted:
* D395 8 8 D_lateral AREA=2.5E-016    ; (523.5 -2317.001 527.5 -2317)CMOSN395 8 8 D_lateral AREA=2.5E-016    
M393 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M392 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M391 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M390 727 724 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M389 724 8 725 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M388 725 8 724 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M387 724 8 725 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M386 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M385 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M384 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M383 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M382 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M381 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M380 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M379 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M378 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M377 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M376 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M375 12 725 727 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M374 12 725 727 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
* Pins of element D372 are shorted:
* D372 12 12 D_lateral AREA=2.5E-016    ; (504.5 -2377 508.5 -2376.999)CMOSN372 12 12 D_lateral AREA=2.5E-016    
* Pins of element D371 are shorted:
* D371 12 12 D_lateral AREA=2.5E-016    ; (488.5 -2377 492.5 -2376.999)CMOSN371 12 12 D_lateral AREA=2.5E-016    
* Pins of element D370 are shorted:
* D370 12 12 D_lateral AREA=2.5E-016    ; (472.5 -2377 476.5 -2376.999)CMOSN370 12 12 D_lateral AREA=2.5E-016    
* Pins of element D369 are shorted:
* D369 12 12 D_lateral AREA=2.5E-016    ; (456.5 -2377 460.5 -2376.999)CMOSN369 12 12 D_lateral AREA=2.5E-016    
* Pins of element D368 are shorted:
* D368 12 12 D_lateral AREA=2.5E-016    ; (440.5 -2377 444.5 -2376.999)CMOSN368 12 12 D_lateral AREA=2.5E-016    
* Pins of element D367 are shorted:
* D367 12 12 D_lateral AREA=2.5E-016    ; (424.5 -2377 428.5 -2376.999)CMOSN367 12 12 D_lateral AREA=2.5E-016    
* Pins of element D365 are shorted:
* D365 8 8 D_lateral AREA=2.5E-016    ; (507.5 -2317.001 511.5 -2317)CMOSN365 8 8 D_lateral AREA=2.5E-016    
* Pins of element D364 are shorted:
* D364 8 8 D_lateral AREA=2.5E-016    ; (491.5 -2317.001 495.5 -2317)CMOSN364 8 8 D_lateral AREA=2.5E-016    
* Pins of element D363 are shorted:
* D363 8 8 D_lateral AREA=1.8125625f    ; (473.499 -2317.001 479.5 -2294)CMOSN363 8 8 D_lateral AREA=1.8125625f    
M362 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M361 725 699 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=4.5p PS=9u    
M360 725 699 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M359 12 699 725 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M358 725 726 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M357 726 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M356 12 727 709 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
M355 709 727 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D354 are shorted:
* D354 12 12 D_lateral AREA=3.75E-016    ; (376.5 -2312.001 382.5 -2312)CMOSN354 12 12 D_lateral AREA=3.75E-016    
* Pins of element D353 are shorted:
* D353 12 12 D_lateral AREA=2f    ; (373.5 -2331 385.5 -2320.999)CMOSN353 12 12 D_lateral AREA=2f    
* Pins of element D352 are shorted:
* D352 12 12 D_lateral AREA=2.4374375f    ; (342.5 -2347 348.5 -2314)CMOSN352 12 12 D_lateral AREA=2.4374375f    
* Pins of element D351 are shorted:
* D351 12 12 D_lateral AREA=2.687375f    ; (326.5 -2349 330.5 -2314)CMOSN351 12 12 D_lateral AREA=2.687375f    
* Pins of element D350 are shorted:
* D350 12 12 D_lateral AREA=2.3749375f    ; (408.5 -2377 412.5 -2343)CMOSN350 12 12 D_lateral AREA=2.3749375f    
* Pins of element D349 are shorted:
* D349 12 12 D_lateral AREA=2.3749375f    ; (318.5 -2350 322.5 -2316)CMOSN349 12 12 D_lateral AREA=2.3749375f    
M348 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M347 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M346 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M345 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M344 708 709 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M343 708 709 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
* Pins of element D342 are shorted:
* D342 12 12 D_lateral AREA=2.5E-016    ; (302.5 -2350 306.5 -2349.999)CMOSN342 12 12 D_lateral AREA=2.5E-016    
* Pins of element D341 are shorted:
* D341 12 12 D_lateral AREA=2.5E-016    ; (286.5 -2350 290.5 -2349.999)CMOSN341 12 12 D_lateral AREA=2.5E-016    
* Pins of element D340 are shorted:
* D340 12 12 D_lateral AREA=2.5E-016    ; (270.5 -2350 274.5 -2349.999)CMOSN340 12 12 D_lateral AREA=2.5E-016    
M339 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M338 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M337 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M336 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M335 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M334 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M333 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M332 710 728 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M331 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M330 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M329 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M328 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M327 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M326 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M325 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M324 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M323 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M322 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M321 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D319 are shorted:
* D319 12 12 D_lateral AREA=3.249875f    ; (100.5 -2377 108.5 -2341)CMOSN319 12 12 D_lateral AREA=3.249875f    
* Pins of element D318 are shorted:
* D318 12 12 D_lateral AREA=2.5E-016    ; (84.5 -2377 88.5 -2376.999)CMOSN318 12 12 D_lateral AREA=2.5E-016    
* Pins of element D317 are shorted:
* D317 12 12 D_lateral AREA=2.5E-016    ; (68.5 -2377 72.5 -2376.999)CMOSN317 12 12 D_lateral AREA=2.5E-016    
* Pins of element D316 are shorted:
* D316 12 12 D_lateral AREA=2.5E-016    ; (52.5 -2377 56.5 -2376.999)CMOSN316 12 12 D_lateral AREA=2.5E-016    
* Pins of element D315 are shorted:
* D315 12 12 D_lateral AREA=2.5E-016    ; (36.5 -2377 40.5 -2376.999)CMOSN315 12 12 D_lateral AREA=2.5E-016    
* Pins of element D314 are shorted:
* D314 12 12 D_lateral AREA=2.5E-016    ; (20.5 -2377 24.5 -2376.999)CMOSN314 12 12 D_lateral AREA=2.5E-016    
* Pins of element D313 are shorted:
* D313 8 8 D_lateral AREA=8.875125f    ; (103.5 -2317.001 107.501 -2181.999)CMOSN313 8 8 D_lateral AREA=8.875125f    
* Pins of element D312 are shorted:
* D312 8 8 D_lateral AREA=2.5E-016    ; (87.5 -2317.001 91.5 -2317)CMOSN312 8 8 D_lateral AREA=2.5E-016    
* Pins of element D311 are shorted:
* D311 8 8 D_lateral AREA=2.5E-016    ; (71.5 -2317.001 75.5 -2317)CMOSN311 8 8 D_lateral AREA=2.5E-016    
* Pins of element D310 are shorted:
* D310 8 8 D_lateral AREA=2.5E-016    ; (55.5 -2317.001 59.5 -2317)CMOSN310 8 8 D_lateral AREA=2.5E-016    
* Pins of element D309 are shorted:
* D309 8 8 D_lateral AREA=1.8125625f    ; (37.499 -2317.001 43.5 -2294)CMOSN309 8 8 D_lateral AREA=1.8125625f    
M308 728 8 729 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M307 729 8 728 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M306 728 8 729 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M305 12 729 710 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M304 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M303 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M302 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M301 710 729 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M300 12 687 729 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M299 729 687 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M298 12 687 729 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M297 729 730 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M296 730 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
* Pins of element D295 are shorted:
* D295 12 12 D_lateral AREA=3.75E-016    ; (-59.5 -2312.001 -53.5 -2312)CMOSN295 12 12 D_lateral AREA=3.75E-016    
* Pins of element D294 are shorted:
* D294 12 12 D_lateral AREA=2f    ; (-62.5 -2331 -50.5 -2320.999)CMOSN294 12 12 D_lateral AREA=2f    
* Pins of element D292 are shorted:
* D292 12 12 D_lateral AREA=2.5E-016    ; (4.5 -2377 8.5 -2376.999)CMOSN292 12 12 D_lateral AREA=2.5E-016    
* Pins of element D291 are shorted:
* D291 12 12 D_lateral AREA=2.5E-016    ; (-11.5 -2377 -7.5 -2376.999)CMOSN291 12 12 D_lateral AREA=2.5E-016    
* Pins of element D290 are shorted:
* D290 12 12 D_lateral AREA=2.3749375f    ; (-27.5 -2377 -23.5 -2343)CMOSN290 12 12 D_lateral AREA=2.3749375f    
M289 12 731 732 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M288 732 731 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M287 12 731 732 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M286 732 731 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M285 12 731 732 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M284 732 731 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M283 12 731 732 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M282 731 710 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=14.3125p PS=20u    
M281 731 710 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D280 are shorted:
* D280 12 12 D_lateral AREA=2.4374375f    ; (-93.5 -2347 -87.5 -2314)CMOSN280 12 12 D_lateral AREA=2.4374375f    
* Pins of element D279 are shorted:
* D279 12 12 D_lateral AREA=2.687375f    ; (-109.5 -2349 -105.5 -2314)CMOSN279 12 12 D_lateral AREA=2.687375f    
* Pins of element D278 are shorted:
* D278 12 12 D_lateral AREA=2.3749375f    ; (-117.5 -2350 -113.5 -2316)CMOSN278 12 12 D_lateral AREA=2.3749375f    
* Pins of element D277 are shorted:
* D277 12 12 D_lateral AREA=2.5E-016    ; (-133.5 -2350 -129.5 -2349.999)CMOSN277 12 12 D_lateral AREA=2.5E-016    
* Pins of element D276 are shorted:
* D276 12 12 D_lateral AREA=2.5E-016    ; (-149.5 -2350 -145.5 -2349.999)CMOSN276 12 12 D_lateral AREA=2.5E-016    
* Pins of element D275 are shorted:
* D275 12 12 D_lateral AREA=2.5E-016    ; (-165.5 -2350 -161.5 -2349.999)CMOSN275 12 12 D_lateral AREA=2.5E-016    
M274 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M273 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M272 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M271 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M270 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M269 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M268 8 733 711 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M267 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M266 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M265 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M264 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M263 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M262 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M261 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D260 are shorted:
* D260 12 12 D_lateral AREA=3.249875f    ; (-335.5 -2377 -327.5 -2341)CMOSN260 12 12 D_lateral AREA=3.249875f    
* Pins of element D259 are shorted:
* D259 12 12 D_lateral AREA=2.5E-016    ; (-351.5 -2377 -347.5 -2376.999)CMOSN259 12 12 D_lateral AREA=2.5E-016    
* Pins of element D258 are shorted:
* D258 12 12 D_lateral AREA=2.5E-016    ; (-367.5 -2377 -363.5 -2376.999)CMOSN258 12 12 D_lateral AREA=2.5E-016    
* Pins of element D257 are shorted:
* D257 12 12 D_lateral AREA=2.5E-016    ; (-383.5 -2377 -379.5 -2376.999)CMOSN257 12 12 D_lateral AREA=2.5E-016    
* Pins of element D256 are shorted:
* D256 8 8 D_lateral AREA=8.875125f    ; (-332.5 -2317.001 -328.499 -2181.999)CMOSN256 8 8 D_lateral AREA=8.875125f    
* Pins of element D255 are shorted:
* D255 8 8 D_lateral AREA=2.5E-016    ; (-348.5 -2317.001 -344.5 -2317)CMOSN255 8 8 D_lateral AREA=2.5E-016    
* Pins of element D254 are shorted:
* D254 8 8 D_lateral AREA=2.5E-016    ; (-364.5 -2317.001 -360.5 -2317)CMOSN254 8 8 D_lateral AREA=2.5E-016    
* Pins of element D253 are shorted:
* D253 8 8 D_lateral AREA=2.5E-016    ; (-380.5 -2317.001 -376.5 -2317)CMOSN253 8 8 D_lateral AREA=2.5E-016    
M252 711 733 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M251 733 8 712 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M250 712 8 733 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M249 733 8 712 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M248 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M247 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M246 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M245 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M244 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M243 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M242 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M241 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M240 711 712 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M239 12 734 712 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M238 712 734 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M237 12 734 712 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M236 712 735 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
* Pins of element D234 are shorted:
* D234 12 12 D_lateral AREA=2.5E-016    ; (-399.5 -2377 -395.5 -2376.999)CMOSN234 12 12 D_lateral AREA=2.5E-016    
* Pins of element D233 are shorted:
* D233 12 12 D_lateral AREA=2.5E-016    ; (-415.5 -2377 -411.5 -2376.999)CMOSN233 12 12 D_lateral AREA=2.5E-016    
* Pins of element D232 are shorted:
* D232 12 12 D_lateral AREA=2.5E-016    ; (-431.5 -2377 -427.5 -2376.999)CMOSN232 12 12 D_lateral AREA=2.5E-016    
* Pins of element D231 are shorted:
* D231 12 12 D_lateral AREA=2.5E-016    ; (-447.5 -2377 -443.5 -2376.999)CMOSN231 12 12 D_lateral AREA=2.5E-016    
* Pins of element D230 are shorted:
* D230 12 12 D_lateral AREA=2.3749375f    ; (-463.5 -2377 -459.5 -2343)CMOSN230 12 12 D_lateral AREA=2.3749375f    
* Pins of element D229 are shorted:
* D229 8 8 D_lateral AREA=1.8125625f    ; (-398.501 -2317.001 -392.5 -2294)CMOSN229 8 8 D_lateral AREA=1.8125625f    
M228 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M227 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M226 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M225 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M224 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M223 735 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M222 12 711 713 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
M221 713 711 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D220 are shorted:
* D220 12 12 D_lateral AREA=3.75E-016    ; (-495.5 -2312.001 -489.5 -2312)CMOSN220 12 12 D_lateral AREA=3.75E-016    
* Pins of element D219 are shorted:
* D219 12 12 D_lateral AREA=2f    ; (-498.5 -2331 -486.5 -2320.999)CMOSN219 12 12 D_lateral AREA=2f    
* Pins of element D218 are shorted:
* D218 12 12 D_lateral AREA=2.4374375f    ; (-529.5 -2347 -523.5 -2314)CMOSN218 12 12 D_lateral AREA=2.4374375f    
* Pins of element D217 are shorted:
* D217 12 12 D_lateral AREA=2.687375f    ; (-545.5 -2349 -541.5 -2314)CMOSN217 12 12 D_lateral AREA=2.687375f    
* Pins of element D216 are shorted:
* D216 12 12 D_lateral AREA=2.3749375f    ; (-553.5 -2350 -549.5 -2316)CMOSN216 12 12 D_lateral AREA=2.3749375f    
* Pins of element D215 are shorted:
* D215 12 12 D_lateral AREA=2.5E-016    ; (-569.5 -2350 -565.5 -2349.999)CMOSN215 12 12 D_lateral AREA=2.5E-016    
* Pins of element D214 are shorted:
* D214 12 12 D_lateral AREA=2.5E-016    ; (-585.5 -2350 -581.5 -2349.999)CMOSN214 12 12 D_lateral AREA=2.5E-016    
M213 736 713 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M212 736 713 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
* Pins of element D211 are shorted:
* D211 12 12 D_lateral AREA=2.5E-016    ; (-601.5 -2350 -597.5 -2349.999)CMOSN211 12 12 D_lateral AREA=2.5E-016    
M210 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M209 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M208 8 737 743 8 CMOSP L=500n W=16u AD=12.3125p PD=17.625u AS=12p PS=17.5u    
M207 743 739 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M206 743 739 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D204 are shorted:
* D204 12 12 D_lateral AREA=3.249875f    ; (-771.5 -2377 -763.5 -2341)CMOSN204 12 12 D_lateral AREA=3.249875f    
* Pins of element D203 are shorted:
* D203 12 12 D_lateral AREA=2.5E-016    ; (-787.5 -2377 -783.5 -2376.999)CMOSN203 12 12 D_lateral AREA=2.5E-016    
* Pins of element D202 are shorted:
* D202 8 8 D_lateral AREA=8.875125f    ; (-768.5 -2317.001 -764.499 -2181.999)CMOSN202 8 8 D_lateral AREA=8.875125f    
* Pins of element D201 are shorted:
* D201 8 8 D_lateral AREA=2.5E-016    ; (-784.5 -2317.001 -780.5 -2317)CMOSN201 8 8 D_lateral AREA=2.5E-016    
M200 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M199 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M198 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M197 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M196 743 737 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M195 737 8 739 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M194 739 8 737 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M193 737 8 739 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M192 743 739 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M191 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M190 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M189 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M188 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M187 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M186 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M185 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M184 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M183 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M182 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M181 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M180 12 739 743 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
* Pins of element D179 are shorted:
* D179 12 12 D_lateral AREA=2.5E-016    ; (-803.5 -2377 -799.5 -2376.999)CMOSN179 12 12 D_lateral AREA=2.5E-016    
* Pins of element D178 are shorted:
* D178 12 12 D_lateral AREA=2.5E-016    ; (-819.5 -2377 -815.5 -2376.999)CMOSN178 12 12 D_lateral AREA=2.5E-016    
* Pins of element D177 are shorted:
* D177 12 12 D_lateral AREA=2.5E-016    ; (-835.5 -2377 -831.5 -2376.999)CMOSN177 12 12 D_lateral AREA=2.5E-016    
* Pins of element D176 are shorted:
* D176 12 12 D_lateral AREA=2.5E-016    ; (-851.5 -2377 -847.5 -2376.999)CMOSN176 12 12 D_lateral AREA=2.5E-016    
* Pins of element D175 are shorted:
* D175 12 12 D_lateral AREA=2.5E-016    ; (-867.5 -2377 -863.5 -2376.999)CMOSN175 12 12 D_lateral AREA=2.5E-016    
* Pins of element D174 are shorted:
* D174 12 12 D_lateral AREA=2.5E-016    ; (-883.5 -2377 -879.5 -2376.999)CMOSN174 12 12 D_lateral AREA=2.5E-016    
* Pins of element D173 are shorted:
* D173 8 8 D_lateral AREA=2.5E-016    ; (-800.5 -2317.001 -796.5 -2317)CMOSN173 8 8 D_lateral AREA=2.5E-016    
* Pins of element D172 are shorted:
* D172 8 8 D_lateral AREA=2.5E-016    ; (-816.5 -2317.001 -812.5 -2317)CMOSN172 8 8 D_lateral AREA=2.5E-016    
* Pins of element D171 are shorted:
* D171 8 8 D_lateral AREA=1.8125625f    ; (-834.501 -2317.001 -828.5 -2294)CMOSN171 8 8 D_lateral AREA=1.8125625f    
M170 743 739 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M169 12 741 739 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M168 739 741 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M167 12 741 739 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M166 739 740 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M165 740 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
M164 12 743 738 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
M163 738 743 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D162 are shorted:
* D162 12 12 D_lateral AREA=3.75E-016    ; (-931.5 -2312.001 -925.5 -2312)CMOSN162 12 12 D_lateral AREA=3.75E-016    
* Pins of element D161 are shorted:
* D161 12 12 D_lateral AREA=2f    ; (-934.5 -2331 -922.5 -2320.999)CMOSN161 12 12 D_lateral AREA=2f    
* Pins of element D160 are shorted:
* D160 12 12 D_lateral AREA=2.4374375f    ; (-965.5 -2347 -959.5 -2314)CMOSN160 12 12 D_lateral AREA=2.4374375f    
* Pins of element D159 are shorted:
* D159 12 12 D_lateral AREA=2.687375f    ; (-981.5 -2349 -977.5 -2314)CMOSN159 12 12 D_lateral AREA=2.687375f    
* Pins of element D158 are shorted:
* D158 12 12 D_lateral AREA=2.3749375f    ; (-899.5 -2377 -895.5 -2343)CMOSN158 12 12 D_lateral AREA=2.3749375f    
M156 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M155 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M154 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M153 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M152 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M151 742 738 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M150 742 738 12 12 CMOSN L=500n W=8u AD=12p PD=19u AS=6.25p PS=10u    
* Pins of element D149 are shorted:
* D149 12 12 D_lateral AREA=2.3749375f    ; (-989.5 -2350 -985.5 -2316)CMOSN149 12 12 D_lateral AREA=2.3749375f    
* Pins of element D148 are shorted:
* D148 12 12 D_lateral AREA=2.5E-016    ; (-1005.5 -2350 -1001.5 -2349.999)CMOSN148 12 12 D_lateral AREA=2.5E-016    
* Pins of element D147 are shorted:
* D147 12 12 D_lateral AREA=2.5E-016    ; (-1021.5 -2350 -1017.5 -2349.999)CMOSN147 12 12 D_lateral AREA=2.5E-016    
* Pins of element D146 are shorted:
* D146 12 12 D_lateral AREA=2.5E-016    ; (-1037.5 -2350 -1033.5 -2349.999)CMOSN146 12 12 D_lateral AREA=2.5E-016    
M145 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=20.8125p PS=35.25u    
M144 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M143 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M142 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M141 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M140 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M139 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=12.3125p PS=17.625u    
M138 750 744 8 8 CMOSP L=500n W=16u AD=12p PD=17.5u AS=25p PS=35.5u    
M137 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=20p PS=22.5u    
M136 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M135 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M134 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M133 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M132 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M131 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M130 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M129 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M128 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
* Pins of element D126 are shorted:
* D126 12 12 D_lateral AREA=3.249875f    ; (-1207.5 -2377 -1199.5 -2341)CMOSN126 12 12 D_lateral AREA=3.249875f    
* Pins of element D125 are shorted:
* D125 12 12 D_lateral AREA=2.5E-016    ; (-1223.5 -2377 -1219.5 -2376.999)CMOSN125 12 12 D_lateral AREA=2.5E-016    
* Pins of element D124 are shorted:
* D124 12 12 D_lateral AREA=2.5E-016    ; (-1239.5 -2377 -1235.5 -2376.999)CMOSN124 12 12 D_lateral AREA=2.5E-016    
* Pins of element D123 are shorted:
* D123 12 12 D_lateral AREA=2.5E-016    ; (-1255.5 -2377 -1251.5 -2376.999)CMOSN123 12 12 D_lateral AREA=2.5E-016    
* Pins of element D122 are shorted:
* D122 12 12 D_lateral AREA=2.5E-016    ; (-1271.5 -2377 -1267.5 -2376.999)CMOSN122 12 12 D_lateral AREA=2.5E-016    
* Pins of element D121 are shorted:
* D121 12 12 D_lateral AREA=2.5E-016    ; (-1287.5 -2377 -1283.5 -2376.999)CMOSN121 12 12 D_lateral AREA=2.5E-016    
* Pins of element D120 are shorted:
* D120 8 8 D_lateral AREA=8.875125f    ; (-1204.5 -2317.001 -1200.499 -2181.999)CMOSN120 8 8 D_lateral AREA=8.875125f    
* Pins of element D119 are shorted:
* D119 8 8 D_lateral AREA=2.5E-016    ; (-1220.5 -2317.001 -1216.5 -2317)CMOSN119 8 8 D_lateral AREA=2.5E-016    
* Pins of element D118 are shorted:
* D118 8 8 D_lateral AREA=2.5E-016    ; (-1236.5 -2317.001 -1232.5 -2317)CMOSN118 8 8 D_lateral AREA=2.5E-016    
* Pins of element D117 are shorted:
* D117 8 8 D_lateral AREA=2.5E-016    ; (-1252.5 -2317.001 -1248.5 -2317)CMOSN117 8 8 D_lateral AREA=2.5E-016    
* Pins of element D116 are shorted:
* D116 8 8 D_lateral AREA=1.8125625f    ; (-1270.501 -2317.001 -1264.5 -2294)CMOSN116 8 8 D_lateral AREA=1.8125625f    
M115 744 8 745 12 CMOSN L=500n W=3.25u AD=4.875p PD=9.5u AS=2.53125p PS=5u    
M114 745 8 744 12 CMOSN L=500n W=3.5u AD=2.53125p PD=5u AS=2.625p PS=5u    
M113 744 8 745 12 CMOSN L=500n W=3.5u AD=2.625p PD=5u AS=5.25p PS=10u    
M112 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M111 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M110 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M109 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M108 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M107 750 745 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=10.5p PS=19.5u    
M106 12 747 745 12 CMOSN L=500n W=3u AD=4.5p PD=9u AS=2.25p PS=4.5u    
M105 745 747 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M104 12 747 745 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=2.25p PS=4.5u    
M103 745 746 12 12 CMOSN L=500n W=3u AD=2.25p PD=4.5u AS=6.0625p PS=10.75u    
M102 746 8 12 12 CMOSN L=500n W=3.75u AD=5.625p PD=10.5u AS=6.0625p PS=10.75u    
* Pins of element D101 are shorted:
* D101 12 12 D_lateral AREA=3.75E-016    ; (-1367.5 -2312.001 -1361.5 -2312)CMOSN101 12 12 D_lateral AREA=3.75E-016    
* Pins of element D100 are shorted:
* D100 12 12 D_lateral AREA=2f    ; (-1370.5 -2331 -1358.5 -2320.999)CMOSN100 12 12 D_lateral AREA=2f    
* Pins of element D99 are shorted:
* D99 12 12 D_lateral AREA=2.5E-016    ; (-1303.5 -2377 -1299.5 -2376.999)CMOSN99 12 12 D_lateral AREA=2.5E-016    
* Pins of element D98 are shorted:
* D98 12 12 D_lateral AREA=2.5E-016    ; (-1319.5 -2377 -1315.5 -2376.999)CMOSN98 12 12 D_lateral AREA=2.5E-016    
* Pins of element D97 are shorted:
* D97 12 12 D_lateral AREA=2.3749375f    ; (-1335.5 -2377 -1331.5 -2343)CMOSN97 12 12 D_lateral AREA=2.3749375f    
M96 12 748 749 12 CMOSN L=500n W=8u AD=10.5p PD=19.5u AS=6p PS=9.5u    
M95 749 748 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M94 12 748 749 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M93 749 748 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M92 12 748 749 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=6p PS=9.5u    
M91 749 748 12 12 CMOSN L=500n W=8u AD=6p PD=9.5u AS=6.25p PS=10u    
M90 12 748 749 12 CMOSN L=500n W=8u AD=6.25p PD=10u AS=12p PS=19u    
M89 12 750 748 12 CMOSN L=500n W=7.75u AD=14.3125p PD=20u AS=5.8125p PS=9.25u    
M88 748 750 12 12 CMOSN L=500n W=7.75u AD=5.8125p PD=9.25u AS=10.25p PS=20u    
* Pins of element D87 are shorted:
* D87 12 12 D_lateral AREA=2.4374375f    ; (-1401.5 -2347 -1395.5 -2314)CMOSN87 12 12 D_lateral AREA=2.4374375f    
* Pins of element D86 are shorted:
* D86 12 12 D_lateral AREA=2.687375f    ; (-1417.5 -2349 -1413.5 -2314)CMOSN86 12 12 D_lateral AREA=2.687375f    
* Pins of element D85 are shorted:
* D85 12 12 D_lateral AREA=2.3749375f    ; (-1425.5 -2350 -1421.5 -2316)CMOSN85 12 12 D_lateral AREA=2.3749375f    
* Pins of element D84 are shorted:
* D84 12 12 D_lateral AREA=2.5E-016    ; (-1441.5 -2350 -1437.5 -2349.999)CMOSN84 12 12 D_lateral AREA=2.5E-016    
* Pins of element D83 are shorted:
* D83 12 12 D_lateral AREA=2.5E-016    ; (-1457.5 -2350 -1453.5 -2349.999)CMOSN83 12 12 D_lateral AREA=2.5E-016    
* Pins of element D82 are shorted:
* D82 12 12 D_lateral AREA=2.5E-016    ; (-1473.5 -2350 -1469.5 -2349.999)CMOSN82 12 12 D_lateral AREA=2.5E-016    
C24 706 12  184.041f    ; (1133.5 -2802 1419.5 -2516)CMOSN.041f    
C20 723 12  184.041f    ; (697.5 -2802 983.5 -2516)CMOSN.041f    
C16 727 12  184.041f    ; (261.5 -2802 547.5 -2516)CMOSN.041f    
C12 710 12  184.041f    ; (-174.5 -2802 111.5 -2516)CMOSN.041f    
C8 711 12  184.041f    ; (-610.5 -2802 -324.5 -2516)CMOSN.041f    
C4 743 12  184.041f    ; (-1046.5 -2802 -760.5 -2516)CMOSN.041f    
C1 750 12  184.041f    ; (-1482.5 -2802 -1196.5 -2516)CMOSN.041f    

* Total Nodes: 750
* Total Elements: 4422
* Total Number of Shorted Elements not written to the SPICE file: 0
* Output Generation Elapsed Time: 0.125 sec
* Total Extract Elapsed Time: 13.672 sec

* INPUTS 
v1 8 0 5v
v2 12 0 0v

v3 45 0 pulse(0v 5v 50n 0.05n 0.05n 250n 100n)
v4 54 0 0v
v5 248 0 0v
v6 442 0 0v
v7 696 0 0v

v8 73 0 5v
v9 83 0 5v
v10 18 0 5v
v11 334 0 5v
v12 37 0 5v
v13 40 0 5v
v14 41 0 pulse(0v 5v 50n 0.05n 0.05n 250n 100n)


* OUTPUTS 
* OUTPUT can be put in trace in simulation 
* 
.op
.tran 0.1ns 200ns
.probe
.END